`timescale 1ns / 1ps

module tb_uart;

    // 1. Khai b�o tham s?
    parameter DATA_WIDTH = 8;
    
    // Clock 50MHz, Baud 115200 -> Prescale = 54
    reg clk = 0;
    reg rst = 0;
    reg [15:0] prescale = 16'd54; 

    // 2. D�y n?i cho User Interface (G?i v�o FIFO TX)
    reg [DATA_WIDTH-1:0] tx_data_in = 0;   // T�n m?i
    reg                  tx_valid_in = 0;  // T�n m?i
    wire                 tx_ready_out;     // T�n m?i

    // 3. D�y n?i cho User Interface (Nh?n t? FIFO RX)
    wire [DATA_WIDTH-1:0] rx_data_out;     // T�n m?i
    wire                  rx_valid_out;    // T�n m?i
    reg                   rx_ready_in = 1; // Lu�n s?n s�ng nh?n

    // 4. D�y v?t l� UART
    wire txd;
    wire rxd;

    // --- SETUP CLOCK 50MHz ---
    always #10 clk = ~clk;

    // --- LOOPBACK: N?i m?m TX v�o tai RX ---
    assign rxd = txd; 

    // --- G?I MODULE UART_FIFO RA CHI?N ---
    // (L?u �: T�n module ph?i tr�ng v?i t�n trong file uart_fifo.v)
    uart_fifo #(
        .DATA_WIDTH(DATA_WIDTH)
    ) uut (
        .clk(clk),
        .rst(rst),
        
        // N?i d�y ph�a G?i (User -> TX FIFO)
        .tx_data_in(tx_data_in),
        .tx_valid_in(tx_valid_in),
        .tx_ready_out(tx_ready_out),
        
        // N?i d�y ph�a Nh?n (RX FIFO -> User)
        .rx_data_out(rx_data_out),
        .rx_valid_out(rx_valid_out),
        .rx_ready_in(rx_ready_in),
        
        // V?t l�
        .rxd(rxd),
        .txd(txd),
        
        // Config
        .prescale(prescale)
    );

    // --- K?CH B?N TEST: G?I NGUY�N CHU?I "HELLO" ---
    initial begin
        // 1. Reset
        $display("--- BAT DAU SIMULATION ---");
        rst = 1;
        #100;
        rst = 0;
        #100;

        // 2. N?p ??n li�n thanh v�o FIFO (G?i 5 byte li�n t?c)
        // FIFO gi�p n� l�m vi?c n�y c?c nhanh, kh�ng c?n ch? UART g?i xong
        
        // G?i 'H' (0x48)
        wait(tx_ready_out); @(posedge clk);
        tx_data_in = 8'h48; tx_valid_in = 1; 
        
        // G?i 'E' (0x45)
        @(posedge clk); // V� FIFO c�n ch?, c? n�m ti?p v�o lu�n
        tx_data_in = 8'h45;
        
        // G?i 'L' (0x4C)
        @(posedge clk);
        tx_data_in = 8'h4C;
        
        // G?i 'L' (0x4C)
        @(posedge clk);
        tx_data_in = 8'h4C;
        
        // G?i 'O' (0x4F)
        @(posedge clk);
        tx_data_in = 8'h4F;
        
        // Ng?t t�n hi?u n?p
        @(posedge clk);
        tx_valid_in = 0;

        $display("--- Da n?p xong 5 ky tu vao FIFO trong tich tac! ---");

        // 3. B�y gi? ng?i xem UART n� t? l�m vi?c (S�ng s? ch?y r?t d�i)
        // N� m? Wave l�n s? th?y txd nh?y m�a li�n t?c
        
        #500000; // ??i ?? l�u cho 5 k� t? ?i qua (Kho?ng 500us)
        
        $display("--- KET THUC ---");
        $stop;
    end

endmodule