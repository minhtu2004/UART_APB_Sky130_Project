// This is the unpowered netlist.
module uart_apb_wrapper (PCLK,
    PENABLE,
    PREADY,
    PRESETn,
    PSEL,
    PSLVERR,
    PWRITE,
    uart_rx,
    uart_tx,
    PADDR,
    PRDATA,
    PWDATA);
 input PCLK;
 input PENABLE;
 output PREADY;
 input PRESETn;
 input PSEL;
 output PSLVERR;
 input PWRITE;
 input uart_rx;
 output uart_tx;
 input [31:0] PADDR;
 output [31:0] PRDATA;
 input [31:0] PWDATA;

 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net42;
 wire net43;
 wire net67;
 wire net66;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire clknet_0_PCLK;
 wire clknet_2_0__leaf_PCLK;
 wire clknet_2_1__leaf_PCLK;
 wire clknet_2_2__leaf_PCLK;
 wire clknet_2_3__leaf_PCLK;
 wire clknet_leaf_0_PCLK;
 wire clknet_leaf_10_PCLK;
 wire clknet_leaf_11_PCLK;
 wire clknet_leaf_12_PCLK;
 wire clknet_leaf_13_PCLK;
 wire clknet_leaf_14_PCLK;
 wire clknet_leaf_15_PCLK;
 wire clknet_leaf_16_PCLK;
 wire clknet_leaf_17_PCLK;
 wire clknet_leaf_18_PCLK;
 wire clknet_leaf_19_PCLK;
 wire clknet_leaf_1_PCLK;
 wire clknet_leaf_20_PCLK;
 wire clknet_leaf_21_PCLK;
 wire clknet_leaf_22_PCLK;
 wire clknet_leaf_23_PCLK;
 wire clknet_leaf_24_PCLK;
 wire clknet_leaf_25_PCLK;
 wire clknet_leaf_26_PCLK;
 wire clknet_leaf_27_PCLK;
 wire clknet_leaf_28_PCLK;
 wire clknet_leaf_29_PCLK;
 wire clknet_leaf_2_PCLK;
 wire clknet_leaf_30_PCLK;
 wire clknet_leaf_31_PCLK;
 wire clknet_leaf_32_PCLK;
 wire clknet_leaf_33_PCLK;
 wire clknet_leaf_34_PCLK;
 wire clknet_leaf_35_PCLK;
 wire clknet_leaf_36_PCLK;
 wire clknet_leaf_3_PCLK;
 wire clknet_leaf_4_PCLK;
 wire clknet_leaf_5_PCLK;
 wire clknet_leaf_6_PCLK;
 wire clknet_leaf_7_PCLK;
 wire clknet_leaf_8_PCLK;
 wire clknet_leaf_9_PCLK;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net5;
 wire net6;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \uart_inst.fifo_rx_inst.mem[0][0] ;
 wire \uart_inst.fifo_rx_inst.mem[0][1] ;
 wire \uart_inst.fifo_rx_inst.mem[0][2] ;
 wire \uart_inst.fifo_rx_inst.mem[0][3] ;
 wire \uart_inst.fifo_rx_inst.mem[0][4] ;
 wire \uart_inst.fifo_rx_inst.mem[0][5] ;
 wire \uart_inst.fifo_rx_inst.mem[0][6] ;
 wire \uart_inst.fifo_rx_inst.mem[0][7] ;
 wire \uart_inst.fifo_rx_inst.mem[10][0] ;
 wire \uart_inst.fifo_rx_inst.mem[10][1] ;
 wire \uart_inst.fifo_rx_inst.mem[10][2] ;
 wire \uart_inst.fifo_rx_inst.mem[10][3] ;
 wire \uart_inst.fifo_rx_inst.mem[10][4] ;
 wire \uart_inst.fifo_rx_inst.mem[10][5] ;
 wire \uart_inst.fifo_rx_inst.mem[10][6] ;
 wire \uart_inst.fifo_rx_inst.mem[10][7] ;
 wire \uart_inst.fifo_rx_inst.mem[11][0] ;
 wire \uart_inst.fifo_rx_inst.mem[11][1] ;
 wire \uart_inst.fifo_rx_inst.mem[11][2] ;
 wire \uart_inst.fifo_rx_inst.mem[11][3] ;
 wire \uart_inst.fifo_rx_inst.mem[11][4] ;
 wire \uart_inst.fifo_rx_inst.mem[11][5] ;
 wire \uart_inst.fifo_rx_inst.mem[11][6] ;
 wire \uart_inst.fifo_rx_inst.mem[11][7] ;
 wire \uart_inst.fifo_rx_inst.mem[12][0] ;
 wire \uart_inst.fifo_rx_inst.mem[12][1] ;
 wire \uart_inst.fifo_rx_inst.mem[12][2] ;
 wire \uart_inst.fifo_rx_inst.mem[12][3] ;
 wire \uart_inst.fifo_rx_inst.mem[12][4] ;
 wire \uart_inst.fifo_rx_inst.mem[12][5] ;
 wire \uart_inst.fifo_rx_inst.mem[12][6] ;
 wire \uart_inst.fifo_rx_inst.mem[12][7] ;
 wire \uart_inst.fifo_rx_inst.mem[13][0] ;
 wire \uart_inst.fifo_rx_inst.mem[13][1] ;
 wire \uart_inst.fifo_rx_inst.mem[13][2] ;
 wire \uart_inst.fifo_rx_inst.mem[13][3] ;
 wire \uart_inst.fifo_rx_inst.mem[13][4] ;
 wire \uart_inst.fifo_rx_inst.mem[13][5] ;
 wire \uart_inst.fifo_rx_inst.mem[13][6] ;
 wire \uart_inst.fifo_rx_inst.mem[13][7] ;
 wire \uart_inst.fifo_rx_inst.mem[14][0] ;
 wire \uart_inst.fifo_rx_inst.mem[14][1] ;
 wire \uart_inst.fifo_rx_inst.mem[14][2] ;
 wire \uart_inst.fifo_rx_inst.mem[14][3] ;
 wire \uart_inst.fifo_rx_inst.mem[14][4] ;
 wire \uart_inst.fifo_rx_inst.mem[14][5] ;
 wire \uart_inst.fifo_rx_inst.mem[14][6] ;
 wire \uart_inst.fifo_rx_inst.mem[14][7] ;
 wire \uart_inst.fifo_rx_inst.mem[15][0] ;
 wire \uart_inst.fifo_rx_inst.mem[15][1] ;
 wire \uart_inst.fifo_rx_inst.mem[15][2] ;
 wire \uart_inst.fifo_rx_inst.mem[15][3] ;
 wire \uart_inst.fifo_rx_inst.mem[15][4] ;
 wire \uart_inst.fifo_rx_inst.mem[15][5] ;
 wire \uart_inst.fifo_rx_inst.mem[15][6] ;
 wire \uart_inst.fifo_rx_inst.mem[15][7] ;
 wire \uart_inst.fifo_rx_inst.mem[1][0] ;
 wire \uart_inst.fifo_rx_inst.mem[1][1] ;
 wire \uart_inst.fifo_rx_inst.mem[1][2] ;
 wire \uart_inst.fifo_rx_inst.mem[1][3] ;
 wire \uart_inst.fifo_rx_inst.mem[1][4] ;
 wire \uart_inst.fifo_rx_inst.mem[1][5] ;
 wire \uart_inst.fifo_rx_inst.mem[1][6] ;
 wire \uart_inst.fifo_rx_inst.mem[1][7] ;
 wire \uart_inst.fifo_rx_inst.mem[2][0] ;
 wire \uart_inst.fifo_rx_inst.mem[2][1] ;
 wire \uart_inst.fifo_rx_inst.mem[2][2] ;
 wire \uart_inst.fifo_rx_inst.mem[2][3] ;
 wire \uart_inst.fifo_rx_inst.mem[2][4] ;
 wire \uart_inst.fifo_rx_inst.mem[2][5] ;
 wire \uart_inst.fifo_rx_inst.mem[2][6] ;
 wire \uart_inst.fifo_rx_inst.mem[2][7] ;
 wire \uart_inst.fifo_rx_inst.mem[3][0] ;
 wire \uart_inst.fifo_rx_inst.mem[3][1] ;
 wire \uart_inst.fifo_rx_inst.mem[3][2] ;
 wire \uart_inst.fifo_rx_inst.mem[3][3] ;
 wire \uart_inst.fifo_rx_inst.mem[3][4] ;
 wire \uart_inst.fifo_rx_inst.mem[3][5] ;
 wire \uart_inst.fifo_rx_inst.mem[3][6] ;
 wire \uart_inst.fifo_rx_inst.mem[3][7] ;
 wire \uart_inst.fifo_rx_inst.mem[4][0] ;
 wire \uart_inst.fifo_rx_inst.mem[4][1] ;
 wire \uart_inst.fifo_rx_inst.mem[4][2] ;
 wire \uart_inst.fifo_rx_inst.mem[4][3] ;
 wire \uart_inst.fifo_rx_inst.mem[4][4] ;
 wire \uart_inst.fifo_rx_inst.mem[4][5] ;
 wire \uart_inst.fifo_rx_inst.mem[4][6] ;
 wire \uart_inst.fifo_rx_inst.mem[4][7] ;
 wire \uart_inst.fifo_rx_inst.mem[5][0] ;
 wire \uart_inst.fifo_rx_inst.mem[5][1] ;
 wire \uart_inst.fifo_rx_inst.mem[5][2] ;
 wire \uart_inst.fifo_rx_inst.mem[5][3] ;
 wire \uart_inst.fifo_rx_inst.mem[5][4] ;
 wire \uart_inst.fifo_rx_inst.mem[5][5] ;
 wire \uart_inst.fifo_rx_inst.mem[5][6] ;
 wire \uart_inst.fifo_rx_inst.mem[5][7] ;
 wire \uart_inst.fifo_rx_inst.mem[6][0] ;
 wire \uart_inst.fifo_rx_inst.mem[6][1] ;
 wire \uart_inst.fifo_rx_inst.mem[6][2] ;
 wire \uart_inst.fifo_rx_inst.mem[6][3] ;
 wire \uart_inst.fifo_rx_inst.mem[6][4] ;
 wire \uart_inst.fifo_rx_inst.mem[6][5] ;
 wire \uart_inst.fifo_rx_inst.mem[6][6] ;
 wire \uart_inst.fifo_rx_inst.mem[6][7] ;
 wire \uart_inst.fifo_rx_inst.mem[7][0] ;
 wire \uart_inst.fifo_rx_inst.mem[7][1] ;
 wire \uart_inst.fifo_rx_inst.mem[7][2] ;
 wire \uart_inst.fifo_rx_inst.mem[7][3] ;
 wire \uart_inst.fifo_rx_inst.mem[7][4] ;
 wire \uart_inst.fifo_rx_inst.mem[7][5] ;
 wire \uart_inst.fifo_rx_inst.mem[7][6] ;
 wire \uart_inst.fifo_rx_inst.mem[7][7] ;
 wire \uart_inst.fifo_rx_inst.mem[8][0] ;
 wire \uart_inst.fifo_rx_inst.mem[8][1] ;
 wire \uart_inst.fifo_rx_inst.mem[8][2] ;
 wire \uart_inst.fifo_rx_inst.mem[8][3] ;
 wire \uart_inst.fifo_rx_inst.mem[8][4] ;
 wire \uart_inst.fifo_rx_inst.mem[8][5] ;
 wire \uart_inst.fifo_rx_inst.mem[8][6] ;
 wire \uart_inst.fifo_rx_inst.mem[8][7] ;
 wire \uart_inst.fifo_rx_inst.mem[9][0] ;
 wire \uart_inst.fifo_rx_inst.mem[9][1] ;
 wire \uart_inst.fifo_rx_inst.mem[9][2] ;
 wire \uart_inst.fifo_rx_inst.mem[9][3] ;
 wire \uart_inst.fifo_rx_inst.mem[9][4] ;
 wire \uart_inst.fifo_rx_inst.mem[9][5] ;
 wire \uart_inst.fifo_rx_inst.mem[9][6] ;
 wire \uart_inst.fifo_rx_inst.mem[9][7] ;
 wire \uart_inst.fifo_rx_inst.read_ptr_reg[0] ;
 wire \uart_inst.fifo_rx_inst.read_ptr_reg[1] ;
 wire \uart_inst.fifo_rx_inst.read_ptr_reg[2] ;
 wire \uart_inst.fifo_rx_inst.read_ptr_reg[3] ;
 wire \uart_inst.fifo_rx_inst.read_ptr_reg[4] ;
 wire \uart_inst.fifo_rx_inst.write_ptr_reg[0] ;
 wire \uart_inst.fifo_rx_inst.write_ptr_reg[1] ;
 wire \uart_inst.fifo_rx_inst.write_ptr_reg[2] ;
 wire \uart_inst.fifo_rx_inst.write_ptr_reg[3] ;
 wire \uart_inst.fifo_rx_inst.write_ptr_reg[4] ;
 wire \uart_inst.fifo_tx_inst.mem[0][0] ;
 wire \uart_inst.fifo_tx_inst.mem[0][1] ;
 wire \uart_inst.fifo_tx_inst.mem[0][2] ;
 wire \uart_inst.fifo_tx_inst.mem[0][3] ;
 wire \uart_inst.fifo_tx_inst.mem[0][4] ;
 wire \uart_inst.fifo_tx_inst.mem[0][5] ;
 wire \uart_inst.fifo_tx_inst.mem[0][6] ;
 wire \uart_inst.fifo_tx_inst.mem[0][7] ;
 wire \uart_inst.fifo_tx_inst.mem[10][0] ;
 wire \uart_inst.fifo_tx_inst.mem[10][1] ;
 wire \uart_inst.fifo_tx_inst.mem[10][2] ;
 wire \uart_inst.fifo_tx_inst.mem[10][3] ;
 wire \uart_inst.fifo_tx_inst.mem[10][4] ;
 wire \uart_inst.fifo_tx_inst.mem[10][5] ;
 wire \uart_inst.fifo_tx_inst.mem[10][6] ;
 wire \uart_inst.fifo_tx_inst.mem[10][7] ;
 wire \uart_inst.fifo_tx_inst.mem[11][0] ;
 wire \uart_inst.fifo_tx_inst.mem[11][1] ;
 wire \uart_inst.fifo_tx_inst.mem[11][2] ;
 wire \uart_inst.fifo_tx_inst.mem[11][3] ;
 wire \uart_inst.fifo_tx_inst.mem[11][4] ;
 wire \uart_inst.fifo_tx_inst.mem[11][5] ;
 wire \uart_inst.fifo_tx_inst.mem[11][6] ;
 wire \uart_inst.fifo_tx_inst.mem[11][7] ;
 wire \uart_inst.fifo_tx_inst.mem[12][0] ;
 wire \uart_inst.fifo_tx_inst.mem[12][1] ;
 wire \uart_inst.fifo_tx_inst.mem[12][2] ;
 wire \uart_inst.fifo_tx_inst.mem[12][3] ;
 wire \uart_inst.fifo_tx_inst.mem[12][4] ;
 wire \uart_inst.fifo_tx_inst.mem[12][5] ;
 wire \uart_inst.fifo_tx_inst.mem[12][6] ;
 wire \uart_inst.fifo_tx_inst.mem[12][7] ;
 wire \uart_inst.fifo_tx_inst.mem[13][0] ;
 wire \uart_inst.fifo_tx_inst.mem[13][1] ;
 wire \uart_inst.fifo_tx_inst.mem[13][2] ;
 wire \uart_inst.fifo_tx_inst.mem[13][3] ;
 wire \uart_inst.fifo_tx_inst.mem[13][4] ;
 wire \uart_inst.fifo_tx_inst.mem[13][5] ;
 wire \uart_inst.fifo_tx_inst.mem[13][6] ;
 wire \uart_inst.fifo_tx_inst.mem[13][7] ;
 wire \uart_inst.fifo_tx_inst.mem[14][0] ;
 wire \uart_inst.fifo_tx_inst.mem[14][1] ;
 wire \uart_inst.fifo_tx_inst.mem[14][2] ;
 wire \uart_inst.fifo_tx_inst.mem[14][3] ;
 wire \uart_inst.fifo_tx_inst.mem[14][4] ;
 wire \uart_inst.fifo_tx_inst.mem[14][5] ;
 wire \uart_inst.fifo_tx_inst.mem[14][6] ;
 wire \uart_inst.fifo_tx_inst.mem[14][7] ;
 wire \uart_inst.fifo_tx_inst.mem[15][0] ;
 wire \uart_inst.fifo_tx_inst.mem[15][1] ;
 wire \uart_inst.fifo_tx_inst.mem[15][2] ;
 wire \uart_inst.fifo_tx_inst.mem[15][3] ;
 wire \uart_inst.fifo_tx_inst.mem[15][4] ;
 wire \uart_inst.fifo_tx_inst.mem[15][5] ;
 wire \uart_inst.fifo_tx_inst.mem[15][6] ;
 wire \uart_inst.fifo_tx_inst.mem[15][7] ;
 wire \uart_inst.fifo_tx_inst.mem[1][0] ;
 wire \uart_inst.fifo_tx_inst.mem[1][1] ;
 wire \uart_inst.fifo_tx_inst.mem[1][2] ;
 wire \uart_inst.fifo_tx_inst.mem[1][3] ;
 wire \uart_inst.fifo_tx_inst.mem[1][4] ;
 wire \uart_inst.fifo_tx_inst.mem[1][5] ;
 wire \uart_inst.fifo_tx_inst.mem[1][6] ;
 wire \uart_inst.fifo_tx_inst.mem[1][7] ;
 wire \uart_inst.fifo_tx_inst.mem[2][0] ;
 wire \uart_inst.fifo_tx_inst.mem[2][1] ;
 wire \uart_inst.fifo_tx_inst.mem[2][2] ;
 wire \uart_inst.fifo_tx_inst.mem[2][3] ;
 wire \uart_inst.fifo_tx_inst.mem[2][4] ;
 wire \uart_inst.fifo_tx_inst.mem[2][5] ;
 wire \uart_inst.fifo_tx_inst.mem[2][6] ;
 wire \uart_inst.fifo_tx_inst.mem[2][7] ;
 wire \uart_inst.fifo_tx_inst.mem[3][0] ;
 wire \uart_inst.fifo_tx_inst.mem[3][1] ;
 wire \uart_inst.fifo_tx_inst.mem[3][2] ;
 wire \uart_inst.fifo_tx_inst.mem[3][3] ;
 wire \uart_inst.fifo_tx_inst.mem[3][4] ;
 wire \uart_inst.fifo_tx_inst.mem[3][5] ;
 wire \uart_inst.fifo_tx_inst.mem[3][6] ;
 wire \uart_inst.fifo_tx_inst.mem[3][7] ;
 wire \uart_inst.fifo_tx_inst.mem[4][0] ;
 wire \uart_inst.fifo_tx_inst.mem[4][1] ;
 wire \uart_inst.fifo_tx_inst.mem[4][2] ;
 wire \uart_inst.fifo_tx_inst.mem[4][3] ;
 wire \uart_inst.fifo_tx_inst.mem[4][4] ;
 wire \uart_inst.fifo_tx_inst.mem[4][5] ;
 wire \uart_inst.fifo_tx_inst.mem[4][6] ;
 wire \uart_inst.fifo_tx_inst.mem[4][7] ;
 wire \uart_inst.fifo_tx_inst.mem[5][0] ;
 wire \uart_inst.fifo_tx_inst.mem[5][1] ;
 wire \uart_inst.fifo_tx_inst.mem[5][2] ;
 wire \uart_inst.fifo_tx_inst.mem[5][3] ;
 wire \uart_inst.fifo_tx_inst.mem[5][4] ;
 wire \uart_inst.fifo_tx_inst.mem[5][5] ;
 wire \uart_inst.fifo_tx_inst.mem[5][6] ;
 wire \uart_inst.fifo_tx_inst.mem[5][7] ;
 wire \uart_inst.fifo_tx_inst.mem[6][0] ;
 wire \uart_inst.fifo_tx_inst.mem[6][1] ;
 wire \uart_inst.fifo_tx_inst.mem[6][2] ;
 wire \uart_inst.fifo_tx_inst.mem[6][3] ;
 wire \uart_inst.fifo_tx_inst.mem[6][4] ;
 wire \uart_inst.fifo_tx_inst.mem[6][5] ;
 wire \uart_inst.fifo_tx_inst.mem[6][6] ;
 wire \uart_inst.fifo_tx_inst.mem[6][7] ;
 wire \uart_inst.fifo_tx_inst.mem[7][0] ;
 wire \uart_inst.fifo_tx_inst.mem[7][1] ;
 wire \uart_inst.fifo_tx_inst.mem[7][2] ;
 wire \uart_inst.fifo_tx_inst.mem[7][3] ;
 wire \uart_inst.fifo_tx_inst.mem[7][4] ;
 wire \uart_inst.fifo_tx_inst.mem[7][5] ;
 wire \uart_inst.fifo_tx_inst.mem[7][6] ;
 wire \uart_inst.fifo_tx_inst.mem[7][7] ;
 wire \uart_inst.fifo_tx_inst.mem[8][0] ;
 wire \uart_inst.fifo_tx_inst.mem[8][1] ;
 wire \uart_inst.fifo_tx_inst.mem[8][2] ;
 wire \uart_inst.fifo_tx_inst.mem[8][3] ;
 wire \uart_inst.fifo_tx_inst.mem[8][4] ;
 wire \uart_inst.fifo_tx_inst.mem[8][5] ;
 wire \uart_inst.fifo_tx_inst.mem[8][6] ;
 wire \uart_inst.fifo_tx_inst.mem[8][7] ;
 wire \uart_inst.fifo_tx_inst.mem[9][0] ;
 wire \uart_inst.fifo_tx_inst.mem[9][1] ;
 wire \uart_inst.fifo_tx_inst.mem[9][2] ;
 wire \uart_inst.fifo_tx_inst.mem[9][3] ;
 wire \uart_inst.fifo_tx_inst.mem[9][4] ;
 wire \uart_inst.fifo_tx_inst.mem[9][5] ;
 wire \uart_inst.fifo_tx_inst.mem[9][6] ;
 wire \uart_inst.fifo_tx_inst.mem[9][7] ;
 wire \uart_inst.fifo_tx_inst.read_ptr_reg[0] ;
 wire \uart_inst.fifo_tx_inst.read_ptr_reg[1] ;
 wire \uart_inst.fifo_tx_inst.read_ptr_reg[2] ;
 wire \uart_inst.fifo_tx_inst.read_ptr_reg[3] ;
 wire \uart_inst.fifo_tx_inst.read_ptr_reg[4] ;
 wire \uart_inst.fifo_tx_inst.write_ptr_reg[0] ;
 wire \uart_inst.fifo_tx_inst.write_ptr_reg[1] ;
 wire \uart_inst.fifo_tx_inst.write_ptr_reg[2] ;
 wire \uart_inst.fifo_tx_inst.write_ptr_reg[3] ;
 wire \uart_inst.fifo_tx_inst.write_ptr_reg[4] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[3] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.data_reg[0] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.data_reg[1] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.data_reg[2] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.data_reg[3] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.data_reg[4] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.data_reg[5] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.data_reg[6] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.data_reg[7] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[0] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[1] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[4] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[7] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.m_axis_tvalid_reg ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[0] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[10] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[11] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[12] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[13] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[14] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[15] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[16] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[17] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[18] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[1] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[2] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[3] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[4] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[5] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[6] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[7] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ;
 wire \uart_inst.uart_core_inst.uart_rx_inst.rxd_reg ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[0] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[1] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[2] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[3] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[0] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[1] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[2] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[3] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[4] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[5] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[6] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[7] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.data_reg[8] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[0] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[10] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[13] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[14] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[15] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[16] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[17] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[18] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[2] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[3] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[4] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[5] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[6] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[7] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[8] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[9] ;
 wire \uart_inst.uart_core_inst.uart_tx_inst.s_axis_tready_reg ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net18));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__inv_2 _1184_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[2] ),
    .Y(_0925_));
 sky130_fd_sc_hd__nand2_1 _1185_ (.A(_0925_),
    .B(\uart_inst.fifo_tx_inst.write_ptr_reg[2] ),
    .Y(_0926_));
 sky130_fd_sc_hd__or2b_1 _1186_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[2] ),
    .B_N(\uart_inst.fifo_tx_inst.read_ptr_reg[2] ),
    .X(_0927_));
 sky130_fd_sc_hd__clkbuf_8 _1187_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[0] ),
    .X(_0928_));
 sky130_fd_sc_hd__or2b_1 _1188_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[0] ),
    .B_N(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__or2b_1 _1189_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[0] ),
    .B_N(\uart_inst.fifo_tx_inst.read_ptr_reg[0] ),
    .X(_0930_));
 sky130_fd_sc_hd__and4_2 _1190_ (.A(_0926_),
    .B(_0927_),
    .C(_0929_),
    .D(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__or2b_1 _1191_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[4] ),
    .B_N(\uart_inst.fifo_tx_inst.write_ptr_reg[4] ),
    .X(_0932_));
 sky130_fd_sc_hd__or2b_1 _1192_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[4] ),
    .B_N(\uart_inst.fifo_tx_inst.read_ptr_reg[4] ),
    .X(_0933_));
 sky130_fd_sc_hd__nand2_2 _1193_ (.A(_0932_),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__nor2_4 _1194_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .B(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ),
    .Y(_0935_));
 sky130_fd_sc_hd__and2_2 _1195_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .B(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ),
    .X(_0936_));
 sky130_fd_sc_hd__nor2_4 _1196_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[3] ),
    .B(\uart_inst.fifo_tx_inst.read_ptr_reg[3] ),
    .Y(_0937_));
 sky130_fd_sc_hd__and2_2 _1197_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[3] ),
    .B(\uart_inst.fifo_tx_inst.read_ptr_reg[3] ),
    .X(_0938_));
 sky130_fd_sc_hd__o22a_2 _1198_ (.A1(_0935_),
    .A2(_0936_),
    .B1(_0937_),
    .B2(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__and3_1 _1199_ (.A(_0931_),
    .B(_0934_),
    .C(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__or4b_4 _1200_ (.A(net2),
    .B(net1),
    .C(net4),
    .D_N(net3),
    .X(_0941_));
 sky130_fd_sc_hd__clkinv_4 _1201_ (.A(\uart_inst.fifo_rx_inst.read_ptr_reg[3] ),
    .Y(_0942_));
 sky130_fd_sc_hd__buf_4 _1202_ (.A(\uart_inst.fifo_rx_inst.read_ptr_reg[0] ),
    .X(_0943_));
 sky130_fd_sc_hd__clkbuf_4 _1203_ (.A(\uart_inst.fifo_rx_inst.read_ptr_reg[1] ),
    .X(_0944_));
 sky130_fd_sc_hd__mux4_1 _1204_ (.A0(\uart_inst.fifo_rx_inst.mem[12][0] ),
    .A1(\uart_inst.fifo_rx_inst.mem[13][0] ),
    .A2(\uart_inst.fifo_rx_inst.mem[14][0] ),
    .A3(\uart_inst.fifo_rx_inst.mem[15][0] ),
    .S0(_0943_),
    .S1(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__mux4_1 _1205_ (.A0(\uart_inst.fifo_rx_inst.mem[8][0] ),
    .A1(\uart_inst.fifo_rx_inst.mem[9][0] ),
    .A2(\uart_inst.fifo_rx_inst.mem[10][0] ),
    .A3(\uart_inst.fifo_rx_inst.mem[11][0] ),
    .S0(_0943_),
    .S1(_0944_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_4 _1206_ (.A(\uart_inst.fifo_rx_inst.read_ptr_reg[2] ),
    .X(_0947_));
 sky130_fd_sc_hd__inv_4 _1207_ (.A(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__mux2_1 _1208_ (.A0(_0945_),
    .A1(_0946_),
    .S(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__nor2_1 _1209_ (.A(_0942_),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__clkbuf_4 _1210_ (.A(\uart_inst.fifo_rx_inst.read_ptr_reg[3] ),
    .X(_0951_));
 sky130_fd_sc_hd__mux4_1 _1211_ (.A0(\uart_inst.fifo_rx_inst.mem[4][0] ),
    .A1(\uart_inst.fifo_rx_inst.mem[5][0] ),
    .A2(\uart_inst.fifo_rx_inst.mem[6][0] ),
    .A3(\uart_inst.fifo_rx_inst.mem[7][0] ),
    .S0(_0943_),
    .S1(_0944_),
    .X(_0952_));
 sky130_fd_sc_hd__mux4_1 _1212_ (.A0(\uart_inst.fifo_rx_inst.mem[0][0] ),
    .A1(\uart_inst.fifo_rx_inst.mem[1][0] ),
    .A2(\uart_inst.fifo_rx_inst.mem[2][0] ),
    .A3(\uart_inst.fifo_rx_inst.mem[3][0] ),
    .S0(_0943_),
    .S1(_0944_),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _1213_ (.A0(_0952_),
    .A1(_0953_),
    .S(_0948_),
    .X(_0954_));
 sky130_fd_sc_hd__nor4_1 _1214_ (.A(net2),
    .B(net1),
    .C(net4),
    .D(net3),
    .Y(_0955_));
 sky130_fd_sc_hd__o21ai_1 _1215_ (.A1(_0951_),
    .A2(_0954_),
    .B1(net41),
    .Y(_0956_));
 sky130_fd_sc_hd__o22ai_4 _1216_ (.A1(_0940_),
    .A2(_0941_),
    .B1(_0950_),
    .B2(_0956_),
    .Y(net18));
 sky130_fd_sc_hd__mux4_1 _1217_ (.A0(\uart_inst.fifo_rx_inst.mem[12][1] ),
    .A1(\uart_inst.fifo_rx_inst.mem[13][1] ),
    .A2(\uart_inst.fifo_rx_inst.mem[14][1] ),
    .A3(\uart_inst.fifo_rx_inst.mem[15][1] ),
    .S0(_0943_),
    .S1(_0944_),
    .X(_0957_));
 sky130_fd_sc_hd__mux4_1 _1218_ (.A0(\uart_inst.fifo_rx_inst.mem[8][1] ),
    .A1(\uart_inst.fifo_rx_inst.mem[9][1] ),
    .A2(\uart_inst.fifo_rx_inst.mem[10][1] ),
    .A3(\uart_inst.fifo_rx_inst.mem[11][1] ),
    .S0(_0943_),
    .S1(_0944_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _1219_ (.A0(_0957_),
    .A1(_0958_),
    .S(_0948_),
    .X(_0959_));
 sky130_fd_sc_hd__clkbuf_4 _1220_ (.A(_0948_),
    .X(_0960_));
 sky130_fd_sc_hd__buf_4 _1221_ (.A(_0943_),
    .X(_0961_));
 sky130_fd_sc_hd__buf_4 _1222_ (.A(_0944_),
    .X(_0962_));
 sky130_fd_sc_hd__mux4_1 _1223_ (.A0(\uart_inst.fifo_rx_inst.mem[4][1] ),
    .A1(\uart_inst.fifo_rx_inst.mem[5][1] ),
    .A2(\uart_inst.fifo_rx_inst.mem[6][1] ),
    .A3(\uart_inst.fifo_rx_inst.mem[7][1] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__nor2_1 _1224_ (.A(_0960_),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__mux4_1 _1225_ (.A0(\uart_inst.fifo_rx_inst.mem[0][1] ),
    .A1(\uart_inst.fifo_rx_inst.mem[1][1] ),
    .A2(\uart_inst.fifo_rx_inst.mem[2][1] ),
    .A3(\uart_inst.fifo_rx_inst.mem[3][1] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_0965_));
 sky130_fd_sc_hd__o21ai_1 _1226_ (.A1(_0947_),
    .A2(_0965_),
    .B1(_0942_),
    .Y(_0966_));
 sky130_fd_sc_hd__o2bb2ai_1 _1227_ (.A1_N(_0951_),
    .A2_N(_0959_),
    .B1(_0964_),
    .B2(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__nor2_2 _1228_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[4] ),
    .B(\uart_inst.fifo_rx_inst.read_ptr_reg[4] ),
    .Y(_0968_));
 sky130_fd_sc_hd__and2_2 _1229_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[4] ),
    .B(\uart_inst.fifo_rx_inst.read_ptr_reg[4] ),
    .X(_0969_));
 sky130_fd_sc_hd__nor2_2 _1230_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[0] ),
    .B(_0943_),
    .Y(_0970_));
 sky130_fd_sc_hd__and2_2 _1231_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[0] ),
    .B(\uart_inst.fifo_rx_inst.read_ptr_reg[0] ),
    .X(_0971_));
 sky130_fd_sc_hd__clkbuf_4 _1232_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[1] ),
    .X(_0972_));
 sky130_fd_sc_hd__nor2_2 _1233_ (.A(_0972_),
    .B(_0944_),
    .Y(_0973_));
 sky130_fd_sc_hd__and2_1 _1234_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[1] ),
    .B(\uart_inst.fifo_rx_inst.read_ptr_reg[1] ),
    .X(_0974_));
 sky130_fd_sc_hd__o22a_4 _1235_ (.A1(_0970_),
    .A2(_0971_),
    .B1(_0973_),
    .B2(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__nor2_1 _1236_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[2] ),
    .B(\uart_inst.fifo_rx_inst.read_ptr_reg[2] ),
    .Y(_0976_));
 sky130_fd_sc_hd__and2_1 _1237_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[2] ),
    .B(\uart_inst.fifo_rx_inst.read_ptr_reg[2] ),
    .X(_0977_));
 sky130_fd_sc_hd__nor2_1 _1238_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .B(\uart_inst.fifo_rx_inst.read_ptr_reg[3] ),
    .Y(_0978_));
 sky130_fd_sc_hd__and2_1 _1239_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .B(\uart_inst.fifo_rx_inst.read_ptr_reg[3] ),
    .X(_0979_));
 sky130_fd_sc_hd__o22a_4 _1240_ (.A1(_0976_),
    .A2(_0977_),
    .B1(_0978_),
    .B2(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__o211ai_4 _1241_ (.A1(_0968_),
    .A2(_0969_),
    .B1(_0975_),
    .C1(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_2 _1242_ (.A(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__o2bb2ai_2 _1243_ (.A1_N(_0967_),
    .A2_N(net377),
    .B1(_0941_),
    .B2(_0982_),
    .Y(net19));
 sky130_fd_sc_hd__mux4_1 _1244_ (.A0(\uart_inst.fifo_rx_inst.mem[12][2] ),
    .A1(\uart_inst.fifo_rx_inst.mem[13][2] ),
    .A2(\uart_inst.fifo_rx_inst.mem[14][2] ),
    .A3(\uart_inst.fifo_rx_inst.mem[15][2] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_0983_));
 sky130_fd_sc_hd__mux4_1 _1245_ (.A0(\uart_inst.fifo_rx_inst.mem[8][2] ),
    .A1(\uart_inst.fifo_rx_inst.mem[9][2] ),
    .A2(\uart_inst.fifo_rx_inst.mem[10][2] ),
    .A3(\uart_inst.fifo_rx_inst.mem[11][2] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _1246_ (.A0(_0983_),
    .A1(_0984_),
    .S(_0948_),
    .X(_0985_));
 sky130_fd_sc_hd__buf_4 _1247_ (.A(_0943_),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_4 _1248_ (.A(_0944_),
    .X(_0987_));
 sky130_fd_sc_hd__mux4_1 _1249_ (.A0(\uart_inst.fifo_rx_inst.mem[0][2] ),
    .A1(\uart_inst.fifo_rx_inst.mem[1][2] ),
    .A2(\uart_inst.fifo_rx_inst.mem[2][2] ),
    .A3(\uart_inst.fifo_rx_inst.mem[3][2] ),
    .S0(_0986_),
    .S1(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__buf_4 _1250_ (.A(_0943_),
    .X(_0989_));
 sky130_fd_sc_hd__buf_4 _1251_ (.A(_0944_),
    .X(_0990_));
 sky130_fd_sc_hd__mux4_1 _1252_ (.A0(\uart_inst.fifo_rx_inst.mem[4][2] ),
    .A1(\uart_inst.fifo_rx_inst.mem[5][2] ),
    .A2(\uart_inst.fifo_rx_inst.mem[6][2] ),
    .A3(\uart_inst.fifo_rx_inst.mem[7][2] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__a21o_1 _1253_ (.A1(_0947_),
    .A2(_0991_),
    .B1(_0951_),
    .X(_0992_));
 sky130_fd_sc_hd__a21o_1 _1254_ (.A1(_0960_),
    .A2(_0988_),
    .B1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__o211a_1 _1255_ (.A1(_0942_),
    .A2(_0985_),
    .B1(net41),
    .C1(_0993_),
    .X(net20));
 sky130_fd_sc_hd__mux4_1 _1256_ (.A0(\uart_inst.fifo_rx_inst.mem[12][3] ),
    .A1(\uart_inst.fifo_rx_inst.mem[13][3] ),
    .A2(\uart_inst.fifo_rx_inst.mem[14][3] ),
    .A3(\uart_inst.fifo_rx_inst.mem[15][3] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_0994_));
 sky130_fd_sc_hd__mux4_1 _1257_ (.A0(\uart_inst.fifo_rx_inst.mem[8][3] ),
    .A1(\uart_inst.fifo_rx_inst.mem[9][3] ),
    .A2(\uart_inst.fifo_rx_inst.mem[10][3] ),
    .A3(\uart_inst.fifo_rx_inst.mem[11][3] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_1 _1258_ (.A0(_0994_),
    .A1(_0995_),
    .S(_0948_),
    .X(_0996_));
 sky130_fd_sc_hd__mux4_1 _1259_ (.A0(\uart_inst.fifo_rx_inst.mem[0][3] ),
    .A1(\uart_inst.fifo_rx_inst.mem[1][3] ),
    .A2(\uart_inst.fifo_rx_inst.mem[2][3] ),
    .A3(\uart_inst.fifo_rx_inst.mem[3][3] ),
    .S0(_0986_),
    .S1(_0987_),
    .X(_0997_));
 sky130_fd_sc_hd__mux4_1 _1260_ (.A0(\uart_inst.fifo_rx_inst.mem[4][3] ),
    .A1(\uart_inst.fifo_rx_inst.mem[5][3] ),
    .A2(\uart_inst.fifo_rx_inst.mem[6][3] ),
    .A3(\uart_inst.fifo_rx_inst.mem[7][3] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_0998_));
 sky130_fd_sc_hd__a21o_1 _1261_ (.A1(_0947_),
    .A2(_0998_),
    .B1(_0951_),
    .X(_0999_));
 sky130_fd_sc_hd__a21o_1 _1262_ (.A1(_0960_),
    .A2(_0997_),
    .B1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__o211a_1 _1263_ (.A1(_0942_),
    .A2(_0996_),
    .B1(net40),
    .C1(_1000_),
    .X(net21));
 sky130_fd_sc_hd__mux4_1 _1264_ (.A0(\uart_inst.fifo_rx_inst.mem[12][4] ),
    .A1(\uart_inst.fifo_rx_inst.mem[13][4] ),
    .A2(\uart_inst.fifo_rx_inst.mem[14][4] ),
    .A3(\uart_inst.fifo_rx_inst.mem[15][4] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_1001_));
 sky130_fd_sc_hd__mux4_1 _1265_ (.A0(\uart_inst.fifo_rx_inst.mem[8][4] ),
    .A1(\uart_inst.fifo_rx_inst.mem[9][4] ),
    .A2(\uart_inst.fifo_rx_inst.mem[10][4] ),
    .A3(\uart_inst.fifo_rx_inst.mem[11][4] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _1266_ (.A0(_1001_),
    .A1(_1002_),
    .S(_0948_),
    .X(_1003_));
 sky130_fd_sc_hd__mux4_1 _1267_ (.A0(\uart_inst.fifo_rx_inst.mem[0][4] ),
    .A1(\uart_inst.fifo_rx_inst.mem[1][4] ),
    .A2(\uart_inst.fifo_rx_inst.mem[2][4] ),
    .A3(\uart_inst.fifo_rx_inst.mem[3][4] ),
    .S0(_0986_),
    .S1(_0987_),
    .X(_1004_));
 sky130_fd_sc_hd__mux4_1 _1268_ (.A0(\uart_inst.fifo_rx_inst.mem[4][4] ),
    .A1(\uart_inst.fifo_rx_inst.mem[5][4] ),
    .A2(\uart_inst.fifo_rx_inst.mem[6][4] ),
    .A3(\uart_inst.fifo_rx_inst.mem[7][4] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_1005_));
 sky130_fd_sc_hd__a21o_1 _1269_ (.A1(_0947_),
    .A2(_1005_),
    .B1(_0951_),
    .X(_1006_));
 sky130_fd_sc_hd__a21o_1 _1270_ (.A1(_0960_),
    .A2(_1004_),
    .B1(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__o211a_1 _1271_ (.A1(_0942_),
    .A2(_1003_),
    .B1(net41),
    .C1(_1007_),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 _1272_ (.A0(\uart_inst.fifo_rx_inst.mem[12][5] ),
    .A1(\uart_inst.fifo_rx_inst.mem[13][5] ),
    .A2(\uart_inst.fifo_rx_inst.mem[14][5] ),
    .A3(\uart_inst.fifo_rx_inst.mem[15][5] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_1008_));
 sky130_fd_sc_hd__mux4_1 _1273_ (.A0(\uart_inst.fifo_rx_inst.mem[8][5] ),
    .A1(\uart_inst.fifo_rx_inst.mem[9][5] ),
    .A2(\uart_inst.fifo_rx_inst.mem[10][5] ),
    .A3(\uart_inst.fifo_rx_inst.mem[11][5] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _1274_ (.A0(_1008_),
    .A1(_1009_),
    .S(_0948_),
    .X(_1010_));
 sky130_fd_sc_hd__mux4_1 _1275_ (.A0(\uart_inst.fifo_rx_inst.mem[0][5] ),
    .A1(\uart_inst.fifo_rx_inst.mem[1][5] ),
    .A2(\uart_inst.fifo_rx_inst.mem[2][5] ),
    .A3(\uart_inst.fifo_rx_inst.mem[3][5] ),
    .S0(_0986_),
    .S1(_0987_),
    .X(_1011_));
 sky130_fd_sc_hd__mux4_1 _1276_ (.A0(\uart_inst.fifo_rx_inst.mem[4][5] ),
    .A1(\uart_inst.fifo_rx_inst.mem[5][5] ),
    .A2(\uart_inst.fifo_rx_inst.mem[6][5] ),
    .A3(\uart_inst.fifo_rx_inst.mem[7][5] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_1012_));
 sky130_fd_sc_hd__a21o_1 _1277_ (.A1(_0947_),
    .A2(_1012_),
    .B1(_0951_),
    .X(_1013_));
 sky130_fd_sc_hd__a21o_1 _1278_ (.A1(_0960_),
    .A2(_1011_),
    .B1(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__o211a_1 _1279_ (.A1(_0942_),
    .A2(_1010_),
    .B1(net40),
    .C1(_1014_),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 _1280_ (.A0(\uart_inst.fifo_rx_inst.mem[12][6] ),
    .A1(\uart_inst.fifo_rx_inst.mem[13][6] ),
    .A2(\uart_inst.fifo_rx_inst.mem[14][6] ),
    .A3(\uart_inst.fifo_rx_inst.mem[15][6] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_1015_));
 sky130_fd_sc_hd__mux4_1 _1281_ (.A0(\uart_inst.fifo_rx_inst.mem[8][6] ),
    .A1(\uart_inst.fifo_rx_inst.mem[9][6] ),
    .A2(\uart_inst.fifo_rx_inst.mem[10][6] ),
    .A3(\uart_inst.fifo_rx_inst.mem[11][6] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _1282_ (.A0(_1015_),
    .A1(_1016_),
    .S(_0948_),
    .X(_1017_));
 sky130_fd_sc_hd__mux4_1 _1283_ (.A0(\uart_inst.fifo_rx_inst.mem[0][6] ),
    .A1(\uart_inst.fifo_rx_inst.mem[1][6] ),
    .A2(\uart_inst.fifo_rx_inst.mem[2][6] ),
    .A3(\uart_inst.fifo_rx_inst.mem[3][6] ),
    .S0(_0986_),
    .S1(_0987_),
    .X(_1018_));
 sky130_fd_sc_hd__mux4_1 _1284_ (.A0(\uart_inst.fifo_rx_inst.mem[4][6] ),
    .A1(\uart_inst.fifo_rx_inst.mem[5][6] ),
    .A2(\uart_inst.fifo_rx_inst.mem[6][6] ),
    .A3(\uart_inst.fifo_rx_inst.mem[7][6] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_1019_));
 sky130_fd_sc_hd__a21o_1 _1285_ (.A1(_0947_),
    .A2(_1019_),
    .B1(_0951_),
    .X(_1020_));
 sky130_fd_sc_hd__a21o_1 _1286_ (.A1(_0960_),
    .A2(_1018_),
    .B1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__o211a_1 _1287_ (.A1(_0942_),
    .A2(_1017_),
    .B1(net40),
    .C1(_1021_),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 _1288_ (.A0(\uart_inst.fifo_rx_inst.mem[12][7] ),
    .A1(\uart_inst.fifo_rx_inst.mem[13][7] ),
    .A2(\uart_inst.fifo_rx_inst.mem[14][7] ),
    .A3(\uart_inst.fifo_rx_inst.mem[15][7] ),
    .S0(_0961_),
    .S1(_0962_),
    .X(_1022_));
 sky130_fd_sc_hd__mux4_1 _1289_ (.A0(\uart_inst.fifo_rx_inst.mem[8][7] ),
    .A1(\uart_inst.fifo_rx_inst.mem[9][7] ),
    .A2(\uart_inst.fifo_rx_inst.mem[10][7] ),
    .A3(\uart_inst.fifo_rx_inst.mem[11][7] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_1 _1290_ (.A0(_1022_),
    .A1(_1023_),
    .S(_0948_),
    .X(_1024_));
 sky130_fd_sc_hd__mux4_1 _1291_ (.A0(\uart_inst.fifo_rx_inst.mem[0][7] ),
    .A1(\uart_inst.fifo_rx_inst.mem[1][7] ),
    .A2(\uart_inst.fifo_rx_inst.mem[2][7] ),
    .A3(\uart_inst.fifo_rx_inst.mem[3][7] ),
    .S0(_0986_),
    .S1(_0987_),
    .X(_1025_));
 sky130_fd_sc_hd__mux4_1 _1292_ (.A0(\uart_inst.fifo_rx_inst.mem[4][7] ),
    .A1(\uart_inst.fifo_rx_inst.mem[5][7] ),
    .A2(\uart_inst.fifo_rx_inst.mem[6][7] ),
    .A3(\uart_inst.fifo_rx_inst.mem[7][7] ),
    .S0(_0989_),
    .S1(_0990_),
    .X(_1026_));
 sky130_fd_sc_hd__a21o_1 _1293_ (.A1(_0947_),
    .A2(_1026_),
    .B1(_0951_),
    .X(_1027_));
 sky130_fd_sc_hd__a21o_1 _1294_ (.A1(_0960_),
    .A2(_1025_),
    .B1(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__o211a_1 _1295_ (.A1(_0942_),
    .A2(_1024_),
    .B1(net40),
    .C1(_1028_),
    .X(net25));
 sky130_fd_sc_hd__xnor2_4 _1296_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[4] ),
    .B(\uart_inst.fifo_tx_inst.read_ptr_reg[4] ),
    .Y(_1029_));
 sky130_fd_sc_hd__inv_2 _1297_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[2] ),
    .Y(_1030_));
 sky130_fd_sc_hd__inv_2 _1298_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[1] ),
    .Y(_1031_));
 sky130_fd_sc_hd__inv_2 _1299_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[0] ),
    .Y(_1032_));
 sky130_fd_sc_hd__and4b_1 _1300_ (.A_N(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[3] ),
    .B(_1030_),
    .C(_1031_),
    .D(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__buf_4 _1301_ (.A(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__nand4_4 _1302_ (.A(_1029_),
    .B(_0939_),
    .C(_0931_),
    .D(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__or4_4 _1303_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[3] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[2] ),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[1] ),
    .D(_1032_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_4 _1304_ (.A(net6),
    .X(_1037_));
 sky130_fd_sc_hd__nor4_1 _1305_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[3] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[2] ),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ),
    .D(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[0] ),
    .Y(_1038_));
 sky130_fd_sc_hd__nor4_1 _1306_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[7] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[6] ),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[5] ),
    .D(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[4] ),
    .Y(_1039_));
 sky130_fd_sc_hd__inv_2 _1307_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[18] ),
    .Y(_1040_));
 sky130_fd_sc_hd__nand3_2 _1308_ (.A(net38),
    .B(net37),
    .C(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__or2_2 _1309_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[17] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[16] ),
    .X(_1042_));
 sky130_fd_sc_hd__nor4_1 _1310_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[15] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .D(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[10] ),
    .Y(_1043_));
 sky130_fd_sc_hd__nor2_2 _1311_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[9] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[8] ),
    .Y(_1044_));
 sky130_fd_sc_hd__nor2_2 _1312_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[14] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[13] ),
    .Y(_1045_));
 sky130_fd_sc_hd__nand4b_2 _1313_ (.A_N(_1042_),
    .B(_1043_),
    .C(_1044_),
    .D(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__nor2_2 _1314_ (.A(_1041_),
    .B(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__and4_1 _1315_ (.A(_1035_),
    .B(_1036_),
    .C(_1037_),
    .D(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__buf_2 _1316_ (.A(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_4 _1317_ (.A(_1034_),
    .X(_1050_));
 sky130_fd_sc_hd__clkbuf_4 _1318_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[0] ),
    .X(_1051_));
 sky130_fd_sc_hd__buf_4 _1319_ (.A(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__clkbuf_4 _1320_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_4 _1321_ (.A(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__o21ai_1 _1322_ (.A1(_1052_),
    .A2(\uart_inst.fifo_tx_inst.mem[14][0] ),
    .B1(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__inv_2 _1323_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[0] ),
    .Y(_1056_));
 sky130_fd_sc_hd__clkbuf_4 _1324_ (.A(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__nor2_1 _1325_ (.A(\uart_inst.fifo_tx_inst.mem[15][0] ),
    .B(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__buf_4 _1326_ (.A(_1056_),
    .X(_1059_));
 sky130_fd_sc_hd__clkbuf_4 _1327_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[0] ),
    .X(_1060_));
 sky130_fd_sc_hd__buf_4 _1328_ (.A(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__o21ba_1 _1329_ (.A1(_1061_),
    .A2(\uart_inst.fifo_tx_inst.mem[12][0] ),
    .B1_N(_1053_),
    .X(_1062_));
 sky130_fd_sc_hd__o21ai_1 _1330_ (.A1(_1059_),
    .A2(\uart_inst.fifo_tx_inst.mem[13][0] ),
    .B1(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__buf_4 _1331_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[2] ),
    .X(_1064_));
 sky130_fd_sc_hd__o211ai_2 _1332_ (.A1(_1055_),
    .A2(_1058_),
    .B1(_1063_),
    .C1(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__buf_4 _1333_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[3] ),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_4 _1334_ (.A(_0925_),
    .X(_1067_));
 sky130_fd_sc_hd__o21ba_1 _1335_ (.A1(_1061_),
    .A2(\uart_inst.fifo_tx_inst.mem[8][0] ),
    .B1_N(_1053_),
    .X(_1068_));
 sky130_fd_sc_hd__o21ai_1 _1336_ (.A1(_1059_),
    .A2(\uart_inst.fifo_tx_inst.mem[9][0] ),
    .B1(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__clkbuf_4 _1337_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ),
    .X(_1070_));
 sky130_fd_sc_hd__o21a_1 _1338_ (.A1(_1061_),
    .A2(\uart_inst.fifo_tx_inst.mem[10][0] ),
    .B1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__o21ai_1 _1339_ (.A1(\uart_inst.fifo_tx_inst.mem[11][0] ),
    .A2(_1059_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__nand3_1 _1340_ (.A(_1067_),
    .B(_1069_),
    .C(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__or4_1 _1341_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[3] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[2] ),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[1] ),
    .D(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[0] ),
    .X(_1074_));
 sky130_fd_sc_hd__buf_4 _1342_ (.A(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__a31oi_2 _1343_ (.A1(_1065_),
    .A2(_1066_),
    .A3(_1073_),
    .B1(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__clkbuf_8 _1344_ (.A(_1060_),
    .X(_1077_));
 sky130_fd_sc_hd__mux4_1 _1345_ (.A0(\uart_inst.fifo_tx_inst.mem[0][0] ),
    .A1(\uart_inst.fifo_tx_inst.mem[1][0] ),
    .A2(\uart_inst.fifo_tx_inst.mem[2][0] ),
    .A3(\uart_inst.fifo_tx_inst.mem[3][0] ),
    .S0(_1077_),
    .S1(_1054_),
    .X(_1078_));
 sky130_fd_sc_hd__nor2_1 _1346_ (.A(_1052_),
    .B(\uart_inst.fifo_tx_inst.mem[6][0] ),
    .Y(_1079_));
 sky130_fd_sc_hd__buf_4 _1347_ (.A(_1053_),
    .X(_1080_));
 sky130_fd_sc_hd__o21ai_1 _1348_ (.A1(\uart_inst.fifo_tx_inst.mem[7][0] ),
    .A2(_1059_),
    .B1(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__nor2_1 _1349_ (.A(_1052_),
    .B(\uart_inst.fifo_tx_inst.mem[4][0] ),
    .Y(_1082_));
 sky130_fd_sc_hd__buf_2 _1350_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ),
    .X(_1083_));
 sky130_fd_sc_hd__clkbuf_4 _1351_ (.A(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__o21bai_1 _1352_ (.A1(\uart_inst.fifo_tx_inst.mem[5][0] ),
    .A2(_1057_),
    .B1_N(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__o221ai_1 _1353_ (.A1(_1079_),
    .A2(_1081_),
    .B1(_1082_),
    .B2(_1085_),
    .C1(_1064_),
    .Y(_1086_));
 sky130_fd_sc_hd__clkinv_4 _1354_ (.A(_1066_),
    .Y(_1087_));
 sky130_fd_sc_hd__o211ai_1 _1355_ (.A1(_1064_),
    .A2(_1078_),
    .B1(_1086_),
    .C1(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__a2bb2oi_1 _1356_ (.A1_N(net186),
    .A2_N(_1050_),
    .B1(_1076_),
    .B2(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__nand4_4 _1357_ (.A(_0931_),
    .B(_0933_),
    .C(_0932_),
    .D(_0939_),
    .Y(_1090_));
 sky130_fd_sc_hd__clkbuf_4 _1358_ (.A(_1047_),
    .X(_1091_));
 sky130_fd_sc_hd__nor2_1 _1359_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[15] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ),
    .Y(_1092_));
 sky130_fd_sc_hd__nor2_1 _1360_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[10] ),
    .Y(_1093_));
 sky130_fd_sc_hd__nand4_4 _1361_ (.A(_1092_),
    .B(_1093_),
    .C(_1044_),
    .D(_1045_),
    .Y(_1094_));
 sky130_fd_sc_hd__nor2_2 _1362_ (.A(_1042_),
    .B(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand3b_2 _1363_ (.A_N(_1041_),
    .B(_1036_),
    .C(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__o21ai_2 _1364_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[0] ),
    .A2(_1047_),
    .B1(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__o2111ai_4 _1365_ (.A1(_1090_),
    .A2(_1075_),
    .B1(_1037_),
    .C1(_1091_),
    .D1(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__o22a_1 _1366_ (.A1(net207),
    .A2(_1049_),
    .B1(_1089_),
    .B2(_1098_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_4 _1367_ (.A(_0925_),
    .X(_1099_));
 sky130_fd_sc_hd__mux4_1 _1368_ (.A0(\uart_inst.fifo_tx_inst.mem[12][1] ),
    .A1(\uart_inst.fifo_tx_inst.mem[13][1] ),
    .A2(\uart_inst.fifo_tx_inst.mem[14][1] ),
    .A3(\uart_inst.fifo_tx_inst.mem[15][1] ),
    .S0(_1077_),
    .S1(_1054_),
    .X(_1100_));
 sky130_fd_sc_hd__buf_4 _1369_ (.A(_1060_),
    .X(_1101_));
 sky130_fd_sc_hd__o21ba_1 _1370_ (.A1(_1101_),
    .A2(\uart_inst.fifo_tx_inst.mem[8][1] ),
    .B1_N(_1053_),
    .X(_1102_));
 sky130_fd_sc_hd__o21ai_1 _1371_ (.A1(_1059_),
    .A2(\uart_inst.fifo_tx_inst.mem[9][1] ),
    .B1(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__buf_4 _1372_ (.A(_1056_),
    .X(_1104_));
 sky130_fd_sc_hd__or2_1 _1373_ (.A(_1051_),
    .B(\uart_inst.fifo_tx_inst.mem[10][1] ),
    .X(_1105_));
 sky130_fd_sc_hd__o211ai_1 _1374_ (.A1(_1104_),
    .A2(\uart_inst.fifo_tx_inst.mem[11][1] ),
    .B1(_1054_),
    .C1(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__a31oi_1 _1375_ (.A1(_1099_),
    .A2(_1103_),
    .A3(_1106_),
    .B1(_1087_),
    .Y(_1107_));
 sky130_fd_sc_hd__o21ai_1 _1376_ (.A1(_1099_),
    .A2(_1100_),
    .B1(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__mux4_1 _1377_ (.A0(\uart_inst.fifo_tx_inst.mem[4][1] ),
    .A1(\uart_inst.fifo_tx_inst.mem[5][1] ),
    .A2(\uart_inst.fifo_tx_inst.mem[6][1] ),
    .A3(\uart_inst.fifo_tx_inst.mem[7][1] ),
    .S0(_1077_),
    .S1(_1054_),
    .X(_1109_));
 sky130_fd_sc_hd__nor2_1 _1378_ (.A(_1052_),
    .B(\uart_inst.fifo_tx_inst.mem[0][1] ),
    .Y(_1110_));
 sky130_fd_sc_hd__o21bai_1 _1379_ (.A1(\uart_inst.fifo_tx_inst.mem[1][1] ),
    .A2(_1104_),
    .B1_N(_1070_),
    .Y(_1111_));
 sky130_fd_sc_hd__o21a_1 _1380_ (.A1(_1101_),
    .A2(\uart_inst.fifo_tx_inst.mem[2][1] ),
    .B1(_1070_),
    .X(_1112_));
 sky130_fd_sc_hd__o21ai_1 _1381_ (.A1(\uart_inst.fifo_tx_inst.mem[3][1] ),
    .A2(_1057_),
    .B1(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__o211ai_1 _1382_ (.A1(_1110_),
    .A2(_1111_),
    .B1(_1067_),
    .C1(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__o211ai_1 _1383_ (.A1(_1099_),
    .A2(_1109_),
    .B1(_1114_),
    .C1(_1087_),
    .Y(_1115_));
 sky130_fd_sc_hd__nor2_1 _1384_ (.A(net180),
    .B(_1050_),
    .Y(_1116_));
 sky130_fd_sc_hd__a31oi_1 _1385_ (.A1(_1108_),
    .A2(_1115_),
    .A3(_1050_),
    .B1(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__o22a_1 _1386_ (.A1(net186),
    .A2(_1049_),
    .B1(_1098_),
    .B2(_1117_),
    .X(_0001_));
 sky130_fd_sc_hd__mux4_1 _1387_ (.A0(\uart_inst.fifo_tx_inst.mem[12][2] ),
    .A1(\uart_inst.fifo_tx_inst.mem[13][2] ),
    .A2(\uart_inst.fifo_tx_inst.mem[14][2] ),
    .A3(\uart_inst.fifo_tx_inst.mem[15][2] ),
    .S0(_1077_),
    .S1(_1054_),
    .X(_1118_));
 sky130_fd_sc_hd__o21ba_1 _1388_ (.A1(_1101_),
    .A2(\uart_inst.fifo_tx_inst.mem[8][2] ),
    .B1_N(_1053_),
    .X(_1119_));
 sky130_fd_sc_hd__o21ai_1 _1389_ (.A1(_1059_),
    .A2(\uart_inst.fifo_tx_inst.mem[9][2] ),
    .B1(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__or2_1 _1390_ (.A(_1051_),
    .B(\uart_inst.fifo_tx_inst.mem[10][2] ),
    .X(_1121_));
 sky130_fd_sc_hd__o211ai_1 _1391_ (.A1(_1104_),
    .A2(\uart_inst.fifo_tx_inst.mem[11][2] ),
    .B1(_1054_),
    .C1(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__a31oi_1 _1392_ (.A1(_1067_),
    .A2(_1120_),
    .A3(_1122_),
    .B1(_1087_),
    .Y(_1123_));
 sky130_fd_sc_hd__o21ai_1 _1393_ (.A1(_1099_),
    .A2(_1118_),
    .B1(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__mux4_1 _1394_ (.A0(\uart_inst.fifo_tx_inst.mem[4][2] ),
    .A1(\uart_inst.fifo_tx_inst.mem[5][2] ),
    .A2(\uart_inst.fifo_tx_inst.mem[6][2] ),
    .A3(\uart_inst.fifo_tx_inst.mem[7][2] ),
    .S0(_1101_),
    .S1(_1084_),
    .X(_1125_));
 sky130_fd_sc_hd__nor2_1 _1395_ (.A(_1052_),
    .B(\uart_inst.fifo_tx_inst.mem[2][2] ),
    .Y(_1126_));
 sky130_fd_sc_hd__o21ai_1 _1396_ (.A1(\uart_inst.fifo_tx_inst.mem[3][2] ),
    .A2(_1104_),
    .B1(_1080_),
    .Y(_1127_));
 sky130_fd_sc_hd__o21ba_1 _1397_ (.A1(_1061_),
    .A2(\uart_inst.fifo_tx_inst.mem[0][2] ),
    .B1_N(_1053_),
    .X(_1128_));
 sky130_fd_sc_hd__o21ai_1 _1398_ (.A1(_1059_),
    .A2(\uart_inst.fifo_tx_inst.mem[1][2] ),
    .B1(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__o211ai_1 _1399_ (.A1(_1126_),
    .A2(_1127_),
    .B1(_1129_),
    .C1(_1067_),
    .Y(_1130_));
 sky130_fd_sc_hd__o211ai_1 _1400_ (.A1(_1099_),
    .A2(_1125_),
    .B1(_1130_),
    .C1(_1087_),
    .Y(_1131_));
 sky130_fd_sc_hd__nor2_1 _1401_ (.A(net175),
    .B(_1034_),
    .Y(_1132_));
 sky130_fd_sc_hd__a31oi_1 _1402_ (.A1(_1124_),
    .A2(_1131_),
    .A3(_1050_),
    .B1(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__o22a_1 _1403_ (.A1(net180),
    .A2(_1049_),
    .B1(_1098_),
    .B2(_1133_),
    .X(_0002_));
 sky130_fd_sc_hd__mux4_1 _1404_ (.A0(\uart_inst.fifo_tx_inst.mem[0][3] ),
    .A1(\uart_inst.fifo_tx_inst.mem[1][3] ),
    .A2(\uart_inst.fifo_tx_inst.mem[2][3] ),
    .A3(\uart_inst.fifo_tx_inst.mem[3][3] ),
    .S0(_1077_),
    .S1(_1054_),
    .X(_1134_));
 sky130_fd_sc_hd__nor2_1 _1405_ (.A(_1052_),
    .B(\uart_inst.fifo_tx_inst.mem[4][3] ),
    .Y(_1135_));
 sky130_fd_sc_hd__o21bai_1 _1406_ (.A1(\uart_inst.fifo_tx_inst.mem[5][3] ),
    .A2(_1059_),
    .B1_N(_1070_),
    .Y(_1136_));
 sky130_fd_sc_hd__o21a_1 _1407_ (.A1(_1101_),
    .A2(\uart_inst.fifo_tx_inst.mem[6][3] ),
    .B1(_1070_),
    .X(_1137_));
 sky130_fd_sc_hd__o21ai_1 _1408_ (.A1(\uart_inst.fifo_tx_inst.mem[7][3] ),
    .A2(_1057_),
    .B1(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__o211ai_1 _1409_ (.A1(_1135_),
    .A2(_1136_),
    .B1(_1064_),
    .C1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__o211ai_2 _1410_ (.A1(_1064_),
    .A2(_1134_),
    .B1(_1139_),
    .C1(_1087_),
    .Y(_1140_));
 sky130_fd_sc_hd__mux4_1 _1411_ (.A0(\uart_inst.fifo_tx_inst.mem[12][3] ),
    .A1(\uart_inst.fifo_tx_inst.mem[13][3] ),
    .A2(\uart_inst.fifo_tx_inst.mem[14][3] ),
    .A3(\uart_inst.fifo_tx_inst.mem[15][3] ),
    .S0(_1101_),
    .S1(_1084_),
    .X(_1141_));
 sky130_fd_sc_hd__o21a_1 _1412_ (.A1(_1101_),
    .A2(\uart_inst.fifo_tx_inst.mem[10][3] ),
    .B1(_1070_),
    .X(_1142_));
 sky130_fd_sc_hd__o21ai_1 _1413_ (.A1(\uart_inst.fifo_tx_inst.mem[11][3] ),
    .A2(_1057_),
    .B1(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__o21ba_1 _1414_ (.A1(_1101_),
    .A2(\uart_inst.fifo_tx_inst.mem[8][3] ),
    .B1_N(_1053_),
    .X(_1144_));
 sky130_fd_sc_hd__o21ai_1 _1415_ (.A1(_1057_),
    .A2(\uart_inst.fifo_tx_inst.mem[9][3] ),
    .B1(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__nand3_1 _1416_ (.A(_1099_),
    .B(_1143_),
    .C(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__o211ai_2 _1417_ (.A1(_1099_),
    .A2(_1141_),
    .B1(_1146_),
    .C1(_1066_),
    .Y(_1147_));
 sky130_fd_sc_hd__nor2_1 _1418_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[4] ),
    .B(_1034_),
    .Y(_1148_));
 sky130_fd_sc_hd__a31oi_1 _1419_ (.A1(_1140_),
    .A2(_1147_),
    .A3(_1050_),
    .B1(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__o22a_1 _1420_ (.A1(net175),
    .A2(_1049_),
    .B1(_1098_),
    .B2(_1149_),
    .X(_0003_));
 sky130_fd_sc_hd__and4_1 _1421_ (.A(_1035_),
    .B(_1036_),
    .C(_1037_),
    .D(_1091_),
    .X(_1150_));
 sky130_fd_sc_hd__o21a_1 _1422_ (.A1(_1077_),
    .A2(\uart_inst.fifo_tx_inst.mem[6][4] ),
    .B1(_1084_),
    .X(_1151_));
 sky130_fd_sc_hd__o21ai_1 _1423_ (.A1(\uart_inst.fifo_tx_inst.mem[7][4] ),
    .A2(_1057_),
    .B1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__o21ba_1 _1424_ (.A1(_1077_),
    .A2(\uart_inst.fifo_tx_inst.mem[4][4] ),
    .B1_N(_1070_),
    .X(_1153_));
 sky130_fd_sc_hd__o21ai_1 _1425_ (.A1(_1057_),
    .A2(\uart_inst.fifo_tx_inst.mem[5][4] ),
    .B1(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__clkbuf_4 _1426_ (.A(_1056_),
    .X(_1155_));
 sky130_fd_sc_hd__o21ba_1 _1427_ (.A1(_1060_),
    .A2(\uart_inst.fifo_tx_inst.mem[0][4] ),
    .B1_N(_1083_),
    .X(_1156_));
 sky130_fd_sc_hd__o21ai_1 _1428_ (.A1(_1155_),
    .A2(\uart_inst.fifo_tx_inst.mem[1][4] ),
    .B1(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__o21a_1 _1429_ (.A1(_1051_),
    .A2(\uart_inst.fifo_tx_inst.mem[2][4] ),
    .B1(_1083_),
    .X(_1158_));
 sky130_fd_sc_hd__o21ai_1 _1430_ (.A1(\uart_inst.fifo_tx_inst.mem[3][4] ),
    .A2(_1155_),
    .B1(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__a31o_1 _1431_ (.A1(_1067_),
    .A2(_1157_),
    .A3(_1159_),
    .B1(_1066_),
    .X(_1160_));
 sky130_fd_sc_hd__a31oi_1 _1432_ (.A1(_1064_),
    .A2(_1152_),
    .A3(_1154_),
    .B1(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__or2_1 _1433_ (.A(_1060_),
    .B(\uart_inst.fifo_tx_inst.mem[8][4] ),
    .X(_1162_));
 sky130_fd_sc_hd__o21ai_1 _1434_ (.A1(_1155_),
    .A2(\uart_inst.fifo_tx_inst.mem[9][4] ),
    .B1(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__or2_1 _1435_ (.A(_1060_),
    .B(\uart_inst.fifo_tx_inst.mem[10][4] ),
    .X(_1164_));
 sky130_fd_sc_hd__o211ai_1 _1436_ (.A1(_1155_),
    .A2(\uart_inst.fifo_tx_inst.mem[11][4] ),
    .B1(_1084_),
    .C1(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__o211ai_1 _1437_ (.A1(_1080_),
    .A2(_1163_),
    .B1(_1165_),
    .C1(_1067_),
    .Y(_1166_));
 sky130_fd_sc_hd__nor2_1 _1438_ (.A(_1052_),
    .B(\uart_inst.fifo_tx_inst.mem[12][4] ),
    .Y(_1167_));
 sky130_fd_sc_hd__o21bai_1 _1439_ (.A1(\uart_inst.fifo_tx_inst.mem[13][4] ),
    .A2(_1155_),
    .B1_N(_1070_),
    .Y(_1168_));
 sky130_fd_sc_hd__o21a_1 _1440_ (.A1(_1051_),
    .A2(\uart_inst.fifo_tx_inst.mem[14][4] ),
    .B1(_1083_),
    .X(_1169_));
 sky130_fd_sc_hd__o21ai_1 _1441_ (.A1(\uart_inst.fifo_tx_inst.mem[15][4] ),
    .A2(_1104_),
    .B1(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__o211ai_1 _1442_ (.A1(_1167_),
    .A2(_1168_),
    .B1(_1170_),
    .C1(\uart_inst.fifo_tx_inst.read_ptr_reg[2] ),
    .Y(_1171_));
 sky130_fd_sc_hd__a31o_1 _1443_ (.A1(_1166_),
    .A2(_1171_),
    .A3(_1066_),
    .B1(_1075_),
    .X(_1172_));
 sky130_fd_sc_hd__o22ai_1 _1444_ (.A1(net152),
    .A2(_1050_),
    .B1(_1161_),
    .B2(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__nor2_1 _1445_ (.A(net214),
    .B(_1049_),
    .Y(_1174_));
 sky130_fd_sc_hd__a21oi_1 _1446_ (.A1(_1150_),
    .A2(_1173_),
    .B1(_1174_),
    .Y(_0004_));
 sky130_fd_sc_hd__mux4_1 _1447_ (.A0(\uart_inst.fifo_tx_inst.mem[12][5] ),
    .A1(\uart_inst.fifo_tx_inst.mem[13][5] ),
    .A2(\uart_inst.fifo_tx_inst.mem[14][5] ),
    .A3(\uart_inst.fifo_tx_inst.mem[15][5] ),
    .S0(_1061_),
    .S1(_1084_),
    .X(_1175_));
 sky130_fd_sc_hd__nor2_1 _1448_ (.A(_1052_),
    .B(\uart_inst.fifo_tx_inst.mem[10][5] ),
    .Y(_1176_));
 sky130_fd_sc_hd__o21ai_1 _1449_ (.A1(\uart_inst.fifo_tx_inst.mem[11][5] ),
    .A2(_1155_),
    .B1(_1084_),
    .Y(_1177_));
 sky130_fd_sc_hd__o21ba_1 _1450_ (.A1(_1051_),
    .A2(\uart_inst.fifo_tx_inst.mem[8][5] ),
    .B1_N(_1083_),
    .X(_1178_));
 sky130_fd_sc_hd__o21ai_1 _1451_ (.A1(_1104_),
    .A2(\uart_inst.fifo_tx_inst.mem[9][5] ),
    .B1(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__o211ai_1 _1452_ (.A1(_1176_),
    .A2(_1177_),
    .B1(_1179_),
    .C1(_1067_),
    .Y(_1180_));
 sky130_fd_sc_hd__o211ai_2 _1453_ (.A1(_1099_),
    .A2(_1175_),
    .B1(_1180_),
    .C1(_1066_),
    .Y(_1181_));
 sky130_fd_sc_hd__mux4_1 _1454_ (.A0(\uart_inst.fifo_tx_inst.mem[0][5] ),
    .A1(\uart_inst.fifo_tx_inst.mem[1][5] ),
    .A2(\uart_inst.fifo_tx_inst.mem[2][5] ),
    .A3(\uart_inst.fifo_tx_inst.mem[3][5] ),
    .S0(_1061_),
    .S1(_1084_),
    .X(_1182_));
 sky130_fd_sc_hd__o21ba_1 _1455_ (.A1(_1051_),
    .A2(\uart_inst.fifo_tx_inst.mem[4][5] ),
    .B1_N(_1083_),
    .X(_1183_));
 sky130_fd_sc_hd__o21ai_1 _1456_ (.A1(_1155_),
    .A2(\uart_inst.fifo_tx_inst.mem[5][5] ),
    .B1(_1183_),
    .Y(_0351_));
 sky130_fd_sc_hd__o21a_1 _1457_ (.A1(_1051_),
    .A2(\uart_inst.fifo_tx_inst.mem[6][5] ),
    .B1(_1083_),
    .X(_0352_));
 sky130_fd_sc_hd__o21ai_1 _1458_ (.A1(\uart_inst.fifo_tx_inst.mem[7][5] ),
    .A2(_1155_),
    .B1(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__a31oi_1 _1459_ (.A1(_0351_),
    .A2(_0353_),
    .A3(\uart_inst.fifo_tx_inst.read_ptr_reg[2] ),
    .B1(_1066_),
    .Y(_0354_));
 sky130_fd_sc_hd__o21ai_1 _1460_ (.A1(_1064_),
    .A2(_1182_),
    .B1(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__nor2_1 _1461_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[6] ),
    .B(_1034_),
    .Y(_0356_));
 sky130_fd_sc_hd__a31o_1 _1462_ (.A1(_1181_),
    .A2(_1034_),
    .A3(_0355_),
    .B1(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__nor2_1 _1463_ (.A(net152),
    .B(_1049_),
    .Y(_0358_));
 sky130_fd_sc_hd__a21oi_1 _1464_ (.A1(_1150_),
    .A2(_0357_),
    .B1(_0358_),
    .Y(_0005_));
 sky130_fd_sc_hd__mux4_1 _1465_ (.A0(\uart_inst.fifo_tx_inst.mem[12][6] ),
    .A1(\uart_inst.fifo_tx_inst.mem[13][6] ),
    .A2(\uart_inst.fifo_tx_inst.mem[14][6] ),
    .A3(\uart_inst.fifo_tx_inst.mem[15][6] ),
    .S0(_1077_),
    .S1(_1054_),
    .X(_0359_));
 sky130_fd_sc_hd__o21ba_1 _1466_ (.A1(_1061_),
    .A2(\uart_inst.fifo_tx_inst.mem[8][6] ),
    .B1_N(_1083_),
    .X(_0360_));
 sky130_fd_sc_hd__o21ai_1 _1467_ (.A1(_1104_),
    .A2(\uart_inst.fifo_tx_inst.mem[9][6] ),
    .B1(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__or2_1 _1468_ (.A(_1051_),
    .B(\uart_inst.fifo_tx_inst.mem[10][6] ),
    .X(_0362_));
 sky130_fd_sc_hd__o211ai_1 _1469_ (.A1(_1104_),
    .A2(\uart_inst.fifo_tx_inst.mem[11][6] ),
    .B1(_1054_),
    .C1(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__a31oi_1 _1470_ (.A1(_1067_),
    .A2(_0361_),
    .A3(_0363_),
    .B1(_1087_),
    .Y(_0364_));
 sky130_fd_sc_hd__o21ai_2 _1471_ (.A1(_1099_),
    .A2(_0359_),
    .B1(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__o21ba_1 _1472_ (.A1(_1051_),
    .A2(\uart_inst.fifo_tx_inst.mem[0][6] ),
    .B1_N(_1083_),
    .X(_0366_));
 sky130_fd_sc_hd__o21ai_1 _1473_ (.A1(_1104_),
    .A2(\uart_inst.fifo_tx_inst.mem[1][6] ),
    .B1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__or2_1 _1474_ (.A(_1060_),
    .B(\uart_inst.fifo_tx_inst.mem[2][6] ),
    .X(_0368_));
 sky130_fd_sc_hd__o211ai_1 _1475_ (.A1(_1104_),
    .A2(\uart_inst.fifo_tx_inst.mem[3][6] ),
    .B1(_1084_),
    .C1(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__a31oi_1 _1476_ (.A1(_1067_),
    .A2(_0367_),
    .A3(_0369_),
    .B1(_1066_),
    .Y(_0370_));
 sky130_fd_sc_hd__o21ba_1 _1477_ (.A1(_1101_),
    .A2(\uart_inst.fifo_tx_inst.mem[4][6] ),
    .B1_N(_1053_),
    .X(_0371_));
 sky130_fd_sc_hd__o21ai_1 _1478_ (.A1(_1057_),
    .A2(\uart_inst.fifo_tx_inst.mem[5][6] ),
    .B1(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__o21a_1 _1479_ (.A1(_1061_),
    .A2(\uart_inst.fifo_tx_inst.mem[6][6] ),
    .B1(_1070_),
    .X(_0373_));
 sky130_fd_sc_hd__o21ai_1 _1480_ (.A1(\uart_inst.fifo_tx_inst.mem[7][6] ),
    .A2(_1057_),
    .B1(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand3_1 _1481_ (.A(_0372_),
    .B(_1064_),
    .C(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__a21oi_1 _1482_ (.A1(_0370_),
    .A2(_0375_),
    .B1(_1075_),
    .Y(_0376_));
 sky130_fd_sc_hd__o2bb2ai_1 _1483_ (.A1_N(_0365_),
    .A2_N(_0376_),
    .B1(net149),
    .B2(_1050_),
    .Y(_0377_));
 sky130_fd_sc_hd__nor2_1 _1484_ (.A(net163),
    .B(_1049_),
    .Y(_0378_));
 sky130_fd_sc_hd__a21oi_1 _1485_ (.A1(_1150_),
    .A2(_0377_),
    .B1(_0378_),
    .Y(_0006_));
 sky130_fd_sc_hd__mux4_1 _1486_ (.A0(\uart_inst.fifo_tx_inst.mem[12][7] ),
    .A1(\uart_inst.fifo_tx_inst.mem[13][7] ),
    .A2(\uart_inst.fifo_tx_inst.mem[14][7] ),
    .A3(\uart_inst.fifo_tx_inst.mem[15][7] ),
    .S0(_1101_),
    .S1(_1084_),
    .X(_0379_));
 sky130_fd_sc_hd__o21ba_1 _1487_ (.A1(_1061_),
    .A2(\uart_inst.fifo_tx_inst.mem[8][7] ),
    .B1_N(_1053_),
    .X(_0380_));
 sky130_fd_sc_hd__o21ai_1 _1488_ (.A1(_1059_),
    .A2(\uart_inst.fifo_tx_inst.mem[9][7] ),
    .B1(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__o21a_1 _1489_ (.A1(_1061_),
    .A2(\uart_inst.fifo_tx_inst.mem[10][7] ),
    .B1(_1070_),
    .X(_0382_));
 sky130_fd_sc_hd__o21ai_1 _1490_ (.A1(\uart_inst.fifo_tx_inst.mem[11][7] ),
    .A2(_1059_),
    .B1(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand3_1 _1491_ (.A(_1067_),
    .B(_0381_),
    .C(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__o211ai_2 _1492_ (.A1(_1099_),
    .A2(_0379_),
    .B1(_0384_),
    .C1(_1066_),
    .Y(_0385_));
 sky130_fd_sc_hd__nor2_1 _1493_ (.A(_1077_),
    .B(\uart_inst.fifo_tx_inst.mem[0][7] ),
    .Y(_0386_));
 sky130_fd_sc_hd__o21bai_1 _1494_ (.A1(\uart_inst.fifo_tx_inst.mem[1][7] ),
    .A2(_1056_),
    .B1_N(_1083_),
    .Y(_0387_));
 sky130_fd_sc_hd__o21a_1 _1495_ (.A1(_1060_),
    .A2(\uart_inst.fifo_tx_inst.mem[2][7] ),
    .B1(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ),
    .X(_0388_));
 sky130_fd_sc_hd__o21ai_1 _1496_ (.A1(\uart_inst.fifo_tx_inst.mem[3][7] ),
    .A2(_1155_),
    .B1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__o211a_1 _1497_ (.A1(_0386_),
    .A2(_0387_),
    .B1(_0389_),
    .C1(_0925_),
    .X(_0390_));
 sky130_fd_sc_hd__o21ba_1 _1498_ (.A1(_1060_),
    .A2(\uart_inst.fifo_tx_inst.mem[4][7] ),
    .B1_N(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ),
    .X(_0391_));
 sky130_fd_sc_hd__o21ai_1 _1499_ (.A1(_1155_),
    .A2(\uart_inst.fifo_tx_inst.mem[5][7] ),
    .B1(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__o21a_1 _1500_ (.A1(_1060_),
    .A2(\uart_inst.fifo_tx_inst.mem[6][7] ),
    .B1(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ),
    .X(_0393_));
 sky130_fd_sc_hd__o21ai_1 _1501_ (.A1(\uart_inst.fifo_tx_inst.mem[7][7] ),
    .A2(_1056_),
    .B1(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__a31o_1 _1502_ (.A1(_0392_),
    .A2(\uart_inst.fifo_tx_inst.read_ptr_reg[2] ),
    .A3(_0394_),
    .B1(_1066_),
    .X(_0395_));
 sky130_fd_sc_hd__o21a_1 _1503_ (.A1(_0390_),
    .A2(_0395_),
    .B1(_1034_),
    .X(_0396_));
 sky130_fd_sc_hd__o2bb2ai_1 _1504_ (.A1_N(_0385_),
    .A2_N(_0396_),
    .B1(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[8] ),
    .B2(_1050_),
    .Y(_0397_));
 sky130_fd_sc_hd__nor2_1 _1505_ (.A(net149),
    .B(_1049_),
    .Y(_0398_));
 sky130_fd_sc_hd__a21oi_1 _1506_ (.A1(_1150_),
    .A2(_0397_),
    .B1(_0398_),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_1 _1507_ (.A(net39),
    .B(_1039_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand3b_4 _1508_ (.A_N(_0399_),
    .B(_1095_),
    .C(_1040_),
    .Y(_0400_));
 sky130_fd_sc_hd__o311a_1 _1509_ (.A1(_0400_),
    .A2(_1090_),
    .A3(_1075_),
    .B1(_1097_),
    .C1(_1037_),
    .X(_0241_));
 sky130_fd_sc_hd__o22ai_4 _1510_ (.A1(_0935_),
    .A2(_0936_),
    .B1(_0937_),
    .B2(_0938_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand4_4 _1511_ (.A(_0926_),
    .B(_0927_),
    .C(_0929_),
    .D(_0930_),
    .Y(_0402_));
 sky130_fd_sc_hd__clkbuf_8 _1512_ (.A(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__o311a_1 _1513_ (.A1(_0934_),
    .A2(_0401_),
    .A3(_0403_),
    .B1(_1091_),
    .C1(_1050_),
    .X(_0404_));
 sky130_fd_sc_hd__a22o_1 _1514_ (.A1(net192),
    .A2(_1098_),
    .B1(_0241_),
    .B2(_0404_),
    .X(_0008_));
 sky130_fd_sc_hd__clkbuf_4 _1515_ (.A(net8),
    .X(_0405_));
 sky130_fd_sc_hd__o221ai_4 _1516_ (.A1(_0935_),
    .A2(_0936_),
    .B1(_0937_),
    .B2(_0938_),
    .C1(_0934_),
    .Y(_0406_));
 sky130_fd_sc_hd__buf_8 _1517_ (.A(net35),
    .X(_0407_));
 sky130_fd_sc_hd__and2_1 _1518_ (.A(net5),
    .B(net7),
    .X(_0408_));
 sky130_fd_sc_hd__and3_1 _1519_ (.A(net16),
    .B(net377),
    .C(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__buf_4 _1520_ (.A(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__buf_8 _1521_ (.A(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_4 _1522_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[2] ),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_4 _1523_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[3] ),
    .X(_0413_));
 sky130_fd_sc_hd__or2b_1 _1524_ (.A(_0412_),
    .B_N(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_1 _1525_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__buf_4 _1526_ (.A(_0928_),
    .X(_0416_));
 sky130_fd_sc_hd__o2111ai_4 _1527_ (.A1(_0403_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0415_),
    .D1(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__mux2_1 _1528_ (.A0(_0405_),
    .A1(net316),
    .S(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _1529_ (.A(_0418_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _1530_ (.A(net9),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _1531_ (.A0(_0419_),
    .A1(net323),
    .S(_0417_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _1532_ (.A(_0420_),
    .X(_0010_));
 sky130_fd_sc_hd__clkbuf_4 _1533_ (.A(net10),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _1534_ (.A0(_0421_),
    .A1(net336),
    .S(_0417_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _1535_ (.A(_0422_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_2 _1536_ (.A(net11),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _1537_ (.A0(_0423_),
    .A1(net341),
    .S(_0417_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _1538_ (.A(_0424_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_2 _1539_ (.A(net12),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(_0425_),
    .A1(net319),
    .S(_0417_),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _1541_ (.A(_0426_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _1542_ (.A(net13),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _1543_ (.A0(_0427_),
    .A1(net294),
    .S(_0417_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _1544_ (.A(_0428_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_4 _1545_ (.A(net14),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _1546_ (.A0(_0429_),
    .A1(net348),
    .S(_0417_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _1547_ (.A(_0430_),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_4 _1548_ (.A(net15),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _1549_ (.A0(_0431_),
    .A1(net302),
    .S(_0417_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _1550_ (.A(_0432_),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _1551_ (.A(_0413_),
    .B(\uart_inst.fifo_tx_inst.write_ptr_reg[2] ),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_4 _1552_ (.A(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__nor2b_4 _1553_ (.A(_0928_),
    .B_N(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .Y(_0435_));
 sky130_fd_sc_hd__o2111ai_4 _1554_ (.A1(_0403_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0434_),
    .D1(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__mux2_1 _1555_ (.A0(_0405_),
    .A1(net313),
    .S(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _1556_ (.A(_0437_),
    .X(_0017_));
 sky130_fd_sc_hd__o21a_1 _1557_ (.A1(_0402_),
    .A2(_0406_),
    .B1(_0410_),
    .X(_0438_));
 sky130_fd_sc_hd__buf_4 _1558_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_4 _1559_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_4 _1560_ (.A(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__nand4b_4 _1561_ (.A_N(_0416_),
    .B(_0439_),
    .C(_0434_),
    .D(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__clkbuf_4 _1562_ (.A(_0928_),
    .X(_0443_));
 sky130_fd_sc_hd__buf_2 _1563_ (.A(_0438_),
    .X(_0444_));
 sky130_fd_sc_hd__and4b_1 _1564_ (.A_N(_0443_),
    .B(net9),
    .C(_0444_),
    .D(_0440_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_4 _1565_ (.A(_0434_),
    .X(_0446_));
 sky130_fd_sc_hd__a22o_1 _1566_ (.A1(net170),
    .A2(_0442_),
    .B1(_0445_),
    .B2(_0446_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(_0421_),
    .A1(net315),
    .S(_0436_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _1568_ (.A(_0447_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _1569_ (.A0(_0423_),
    .A1(net335),
    .S(_0436_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _1570_ (.A(_0448_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _1571_ (.A0(_0425_),
    .A1(net297),
    .S(_0436_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _1572_ (.A(_0449_),
    .X(_0021_));
 sky130_fd_sc_hd__o311a_1 _1573_ (.A1(_1029_),
    .A2(_0401_),
    .A3(_0403_),
    .B1(_0411_),
    .C1(_0435_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_4 _1574_ (.A(_0413_),
    .X(_0451_));
 sky130_fd_sc_hd__and3_1 _1575_ (.A(_0451_),
    .B(_0412_),
    .C(net13),
    .X(_0452_));
 sky130_fd_sc_hd__a22o_1 _1576_ (.A1(_0450_),
    .A2(_0452_),
    .B1(_0442_),
    .B2(net159),
    .X(_0022_));
 sky130_fd_sc_hd__and4b_1 _1577_ (.A_N(_0443_),
    .B(net14),
    .C(_0444_),
    .D(_0440_),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _1578_ (.A1(net151),
    .A2(_0442_),
    .B1(_0453_),
    .B2(_0446_),
    .X(_0023_));
 sky130_fd_sc_hd__and4b_1 _1579_ (.A_N(_0443_),
    .B(net15),
    .C(_0444_),
    .D(_0440_),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _1580_ (.A1(net139),
    .A2(_0442_),
    .B1(_0454_),
    .B2(_0446_),
    .X(_0024_));
 sky130_fd_sc_hd__and3b_1 _1581_ (.A_N(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .B(_0412_),
    .C(_0413_),
    .X(_0455_));
 sky130_fd_sc_hd__o2111ai_4 _1582_ (.A1(_0403_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0455_),
    .D1(_0416_),
    .Y(_0456_));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(_0405_),
    .A1(net290),
    .S(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _1584_ (.A(_0457_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1585_ (.A0(_0419_),
    .A1(net287),
    .S(_0456_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _1586_ (.A(_0458_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _1587_ (.A0(_0421_),
    .A1(net279),
    .S(_0456_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _1588_ (.A(_0459_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1589_ (.A0(_0423_),
    .A1(net300),
    .S(_0456_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _1590_ (.A(_0460_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1591_ (.A0(_0425_),
    .A1(net295),
    .S(_0456_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _1592_ (.A(_0461_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1593_ (.A0(_0427_),
    .A1(net325),
    .S(_0456_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _1594_ (.A(_0462_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1595_ (.A0(_0429_),
    .A1(net275),
    .S(_0456_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _1596_ (.A(_0463_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1597_ (.A0(_0431_),
    .A1(net289),
    .S(_0456_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_1 _1598_ (.A(_0464_),
    .X(_0032_));
 sky130_fd_sc_hd__buf_6 _1599_ (.A(_0402_),
    .X(_0465_));
 sky130_fd_sc_hd__nor2_4 _1600_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .B(_0928_),
    .Y(_0466_));
 sky130_fd_sc_hd__o2111ai_4 _1601_ (.A1(_0465_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0434_),
    .D1(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__mux2_1 _1602_ (.A0(_0405_),
    .A1(net312),
    .S(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _1603_ (.A(_0468_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1604_ (.A0(_0419_),
    .A1(net318),
    .S(_0467_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _1605_ (.A(_0469_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(_0421_),
    .A1(net281),
    .S(_0467_),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_1 _1607_ (.A(_0470_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(_0423_),
    .A1(net291),
    .S(_0467_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _1609_ (.A(_0471_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(_0425_),
    .A1(net340),
    .S(_0467_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _1611_ (.A(_0472_),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_4 _1612_ (.A(_0438_),
    .X(_0473_));
 sky130_fd_sc_hd__a32o_1 _1613_ (.A1(_0473_),
    .A2(_0452_),
    .A3(_0466_),
    .B1(_0467_),
    .B2(net154),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _1614_ (.A0(_0429_),
    .A1(net257),
    .S(_0467_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _1615_ (.A(_0474_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(_0431_),
    .A1(net258),
    .S(_0467_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _1617_ (.A(_0475_),
    .X(_0040_));
 sky130_fd_sc_hd__nor2_4 _1618_ (.A(_0968_),
    .B(_0969_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_1 _1619_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[0] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tvalid_reg ),
    .Y(_0477_));
 sky130_fd_sc_hd__a31oi_4 _1620_ (.A1(_0476_),
    .A2(_0975_),
    .A3(_0980_),
    .B1(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__buf_4 _1621_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[2] ),
    .X(_0479_));
 sky130_fd_sc_hd__and3_1 _1622_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .B(_0479_),
    .C(_0972_),
    .X(_0480_));
 sky130_fd_sc_hd__nand2_4 _1623_ (.A(_0478_),
    .B(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__buf_2 _1624_ (.A(_0972_),
    .X(_0482_));
 sky130_fd_sc_hd__buf_2 _1625_ (.A(_0478_),
    .X(_0483_));
 sky130_fd_sc_hd__and3_2 _1626_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[0] ),
    .B(_0482_),
    .C(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__and2_1 _1627_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .B(\uart_inst.fifo_rx_inst.write_ptr_reg[2] ),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_2 _1628_ (.A(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_4 _1629_ (.A(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _1630_ (.A1(net148),
    .A2(_0481_),
    .B1(_0484_),
    .B2(_0487_),
    .X(_0041_));
 sky130_fd_sc_hd__and3_1 _1631_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[1] ),
    .B(_0482_),
    .C(_0483_),
    .X(_0488_));
 sky130_fd_sc_hd__a22o_1 _1632_ (.A1(net166),
    .A2(_0481_),
    .B1(_0488_),
    .B2(_0487_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_4 _1633_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _1634_ (.A0(_0489_),
    .A1(net274),
    .S(_0481_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _1635_ (.A(_0490_),
    .X(_0043_));
 sky130_fd_sc_hd__buf_4 _1636_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _1637_ (.A0(_0491_),
    .A1(net299),
    .S(_0481_),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_1 _1638_ (.A(_0492_),
    .X(_0044_));
 sky130_fd_sc_hd__and3_1 _1639_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[4] ),
    .B(_0482_),
    .C(_0483_),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _1640_ (.A1(net161),
    .A2(_0481_),
    .B1(_0493_),
    .B2(_0487_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_4 _1641_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _1642_ (.A0(_0494_),
    .A1(net314),
    .S(_0481_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _1643_ (.A(_0495_),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_4 _1644_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _1645_ (.A0(_0496_),
    .A1(net283),
    .S(_0481_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_1 _1646_ (.A(_0497_),
    .X(_0047_));
 sky130_fd_sc_hd__and3_1 _1647_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[7] ),
    .B(_0972_),
    .C(_0478_),
    .X(_0498_));
 sky130_fd_sc_hd__a22o_1 _1648_ (.A1(net153),
    .A2(_0481_),
    .B1(_0498_),
    .B2(_0487_),
    .X(_0048_));
 sky130_fd_sc_hd__nor2b_4 _1649_ (.A(_0412_),
    .B_N(_0413_),
    .Y(_0499_));
 sky130_fd_sc_hd__clkbuf_4 _1650_ (.A(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__o2111a_2 _1651_ (.A1(_0465_),
    .A2(_0406_),
    .B1(_0410_),
    .C1(_0928_),
    .D1(_0440_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_4 _1652_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__o2111ai_4 _1653_ (.A1(_0402_),
    .A2(net35),
    .B1(_0410_),
    .C1(_0928_),
    .D1(_0440_),
    .Y(_0503_));
 sky130_fd_sc_hd__clkbuf_4 _1654_ (.A(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__o21a_1 _1655_ (.A1(_0414_),
    .A2(_0504_),
    .B1(net229),
    .X(_0505_));
 sky130_fd_sc_hd__a31o_1 _1656_ (.A1(_0405_),
    .A2(_0500_),
    .A3(_0502_),
    .B1(_0505_),
    .X(_0049_));
 sky130_fd_sc_hd__clkbuf_4 _1657_ (.A(_0440_),
    .X(_0506_));
 sky130_fd_sc_hd__nand4_4 _1658_ (.A(_0506_),
    .B(_0443_),
    .C(_0499_),
    .D(_0439_),
    .Y(_0507_));
 sky130_fd_sc_hd__and4_1 _1659_ (.A(_0506_),
    .B(_0443_),
    .C(net9),
    .D(_0439_),
    .X(_0508_));
 sky130_fd_sc_hd__a22o_1 _1660_ (.A1(net169),
    .A2(_0507_),
    .B1(_0508_),
    .B2(_0500_),
    .X(_0050_));
 sky130_fd_sc_hd__and4_2 _1661_ (.A(_0506_),
    .B(_0416_),
    .C(net10),
    .D(_0444_),
    .X(_0509_));
 sky130_fd_sc_hd__a22o_1 _1662_ (.A1(net171),
    .A2(_0507_),
    .B1(_0509_),
    .B2(_0500_),
    .X(_0051_));
 sky130_fd_sc_hd__o21a_1 _1663_ (.A1(_0414_),
    .A2(_0503_),
    .B1(net241),
    .X(_0510_));
 sky130_fd_sc_hd__a31o_1 _1664_ (.A1(_0423_),
    .A2(_0500_),
    .A3(_0502_),
    .B1(_0510_),
    .X(_0052_));
 sky130_fd_sc_hd__and4_1 _1665_ (.A(_0506_),
    .B(_0443_),
    .C(net12),
    .D(_0439_),
    .X(_0511_));
 sky130_fd_sc_hd__a22o_1 _1666_ (.A1(net206),
    .A2(_0507_),
    .B1(_0511_),
    .B2(_0500_),
    .X(_0053_));
 sky130_fd_sc_hd__and4_1 _1667_ (.A(_0506_),
    .B(_0443_),
    .C(net13),
    .D(_0444_),
    .X(_0512_));
 sky130_fd_sc_hd__a22o_1 _1668_ (.A1(net196),
    .A2(_0507_),
    .B1(_0512_),
    .B2(_0500_),
    .X(_0054_));
 sky130_fd_sc_hd__and4_1 _1669_ (.A(_0506_),
    .B(_0416_),
    .C(net14),
    .D(_0444_),
    .X(_0513_));
 sky130_fd_sc_hd__a22o_1 _1670_ (.A1(net197),
    .A2(_0507_),
    .B1(_0513_),
    .B2(_0500_),
    .X(_0055_));
 sky130_fd_sc_hd__o21a_1 _1671_ (.A1(_0414_),
    .A2(_0503_),
    .B1(net235),
    .X(_0514_));
 sky130_fd_sc_hd__a31o_1 _1672_ (.A1(_0431_),
    .A2(_0500_),
    .A3(_0502_),
    .B1(_0514_),
    .X(_0056_));
 sky130_fd_sc_hd__o2111ai_4 _1673_ (.A1(_0465_),
    .A2(net35),
    .B1(_0499_),
    .C1(_0410_),
    .D1(_0435_),
    .Y(_0515_));
 sky130_fd_sc_hd__mux2_1 _1674_ (.A0(_0405_),
    .A1(net360),
    .S(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _1675_ (.A(_0516_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1676_ (.A0(_0419_),
    .A1(net263),
    .S(_0515_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _1677_ (.A(_0517_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1678_ (.A0(_0421_),
    .A1(net265),
    .S(_0515_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _1679_ (.A(_0518_),
    .X(_0059_));
 sky130_fd_sc_hd__and4b_1 _1680_ (.A_N(_0443_),
    .B(net11),
    .C(_0444_),
    .D(_0440_),
    .X(_0519_));
 sky130_fd_sc_hd__a22o_1 _1681_ (.A1(net189),
    .A2(_0515_),
    .B1(_0519_),
    .B2(_0500_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1682_ (.A0(_0425_),
    .A1(net247),
    .S(_0515_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_1 _1683_ (.A(_0520_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1684_ (.A0(_0427_),
    .A1(net353),
    .S(_0515_),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_1 _1685_ (.A(_0521_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1686_ (.A0(_0429_),
    .A1(net254),
    .S(_0515_),
    .X(_0522_));
 sky130_fd_sc_hd__clkbuf_1 _1687_ (.A(_0522_),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_1 _1688_ (.A1(net173),
    .A2(_0515_),
    .B1(_0454_),
    .B2(_0500_),
    .X(_0064_));
 sky130_fd_sc_hd__nor2_2 _1689_ (.A(_0413_),
    .B(_0412_),
    .Y(_0523_));
 sky130_fd_sc_hd__o2111ai_4 _1690_ (.A1(_0403_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0466_),
    .D1(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__mux2_1 _1691_ (.A0(_0405_),
    .A1(net320),
    .S(net30),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_1 _1692_ (.A(_0525_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1693_ (.A0(_0419_),
    .A1(net350),
    .S(net30),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _1694_ (.A(_0526_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1695_ (.A0(_0421_),
    .A1(net363),
    .S(net30),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _1696_ (.A(_0527_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1697_ (.A0(_0423_),
    .A1(net277),
    .S(net30),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_1 _1698_ (.A(_0528_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1699_ (.A0(_0425_),
    .A1(net349),
    .S(_0524_),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_1 _1700_ (.A(_0529_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1701_ (.A0(_0427_),
    .A1(net324),
    .S(_0524_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_1 _1702_ (.A(_0530_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1703_ (.A0(_0429_),
    .A1(net352),
    .S(_0524_),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_1 _1704_ (.A(_0531_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(_0431_),
    .A1(net307),
    .S(_0524_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _1706_ (.A(_0532_),
    .X(_0072_));
 sky130_fd_sc_hd__o2111ai_4 _1707_ (.A1(_0465_),
    .A2(_0407_),
    .B1(_0499_),
    .C1(_0410_),
    .D1(_0466_),
    .Y(_0533_));
 sky130_fd_sc_hd__mux2_1 _1708_ (.A0(_0405_),
    .A1(net329),
    .S(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_1 _1709_ (.A(_0534_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1710_ (.A0(_0419_),
    .A1(net309),
    .S(_0533_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _1711_ (.A(_0535_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1712_ (.A0(_0421_),
    .A1(net326),
    .S(_0533_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1713_ (.A(_0536_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1714_ (.A0(_0423_),
    .A1(net342),
    .S(_0533_),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_1 _1715_ (.A(_0537_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1716_ (.A0(_0425_),
    .A1(net272),
    .S(net29),
    .X(_0538_));
 sky130_fd_sc_hd__clkbuf_1 _1717_ (.A(_0538_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1718_ (.A0(_0427_),
    .A1(net317),
    .S(net29),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_1 _1719_ (.A(_0539_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1720_ (.A0(_0429_),
    .A1(net346),
    .S(net29),
    .X(_0540_));
 sky130_fd_sc_hd__clkbuf_1 _1721_ (.A(_0540_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1722_ (.A0(_0431_),
    .A1(net301),
    .S(net29),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_1 _1723_ (.A(_0541_),
    .X(_0080_));
 sky130_fd_sc_hd__or2b_1 _1724_ (.A(_0413_),
    .B_N(\uart_inst.fifo_tx_inst.write_ptr_reg[2] ),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_4 _1725_ (.A(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_4 _1726_ (.A(_0416_),
    .X(_0544_));
 sky130_fd_sc_hd__nor2b_4 _1727_ (.A(_0413_),
    .B_N(_0412_),
    .Y(_0545_));
 sky130_fd_sc_hd__clkbuf_4 _1728_ (.A(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__a41o_1 _1729_ (.A1(_0441_),
    .A2(_0544_),
    .A3(_0473_),
    .A4(_0546_),
    .B1(net239),
    .X(_0547_));
 sky130_fd_sc_hd__o31a_1 _1730_ (.A1(_0405_),
    .A2(_0504_),
    .A3(_0543_),
    .B1(_0547_),
    .X(_0081_));
 sky130_fd_sc_hd__a41o_1 _1731_ (.A1(_0441_),
    .A2(_0544_),
    .A3(_0473_),
    .A4(_0546_),
    .B1(net223),
    .X(_0548_));
 sky130_fd_sc_hd__o31a_1 _1732_ (.A1(_0419_),
    .A2(_0504_),
    .A3(_0543_),
    .B1(_0548_),
    .X(_0082_));
 sky130_fd_sc_hd__a41o_1 _1733_ (.A1(_0441_),
    .A2(_0544_),
    .A3(_0473_),
    .A4(_0546_),
    .B1(net224),
    .X(_0549_));
 sky130_fd_sc_hd__o31a_1 _1734_ (.A1(_0421_),
    .A2(_0504_),
    .A3(_0543_),
    .B1(_0549_),
    .X(_0083_));
 sky130_fd_sc_hd__a41o_1 _1735_ (.A1(_0441_),
    .A2(_0544_),
    .A3(_0473_),
    .A4(_0546_),
    .B1(net238),
    .X(_0550_));
 sky130_fd_sc_hd__o31a_1 _1736_ (.A1(_0423_),
    .A2(_0504_),
    .A3(_0543_),
    .B1(_0550_),
    .X(_0084_));
 sky130_fd_sc_hd__a41o_1 _1737_ (.A1(_0441_),
    .A2(_0544_),
    .A3(_0473_),
    .A4(_0546_),
    .B1(net233),
    .X(_0551_));
 sky130_fd_sc_hd__o31a_1 _1738_ (.A1(_0425_),
    .A2(_0504_),
    .A3(_0543_),
    .B1(_0551_),
    .X(_0085_));
 sky130_fd_sc_hd__a41o_1 _1739_ (.A1(_0441_),
    .A2(_0544_),
    .A3(_0439_),
    .A4(_0546_),
    .B1(net248),
    .X(_0552_));
 sky130_fd_sc_hd__o31a_1 _1740_ (.A1(_0427_),
    .A2(_0504_),
    .A3(_0543_),
    .B1(_0552_),
    .X(_0086_));
 sky130_fd_sc_hd__a41o_1 _1741_ (.A1(_0441_),
    .A2(_0544_),
    .A3(_0439_),
    .A4(_0545_),
    .B1(net237),
    .X(_0553_));
 sky130_fd_sc_hd__o31a_1 _1742_ (.A1(_0429_),
    .A2(_0504_),
    .A3(_0543_),
    .B1(_0553_),
    .X(_0087_));
 sky130_fd_sc_hd__a41o_1 _1743_ (.A1(_0441_),
    .A2(_0544_),
    .A3(_0439_),
    .A4(_0545_),
    .B1(net243),
    .X(_0554_));
 sky130_fd_sc_hd__o31a_1 _1744_ (.A1(_0431_),
    .A2(_0504_),
    .A3(_0543_),
    .B1(_0554_),
    .X(_0088_));
 sky130_fd_sc_hd__o2111ai_4 _1745_ (.A1(_0403_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0435_),
    .D1(_0545_),
    .Y(_0555_));
 sky130_fd_sc_hd__mux2_1 _1746_ (.A0(_0405_),
    .A1(net338),
    .S(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__clkbuf_1 _1747_ (.A(_0556_),
    .X(_0089_));
 sky130_fd_sc_hd__nand4b_4 _1748_ (.A_N(_0416_),
    .B(_0439_),
    .C(_0545_),
    .D(_0506_),
    .Y(_0557_));
 sky130_fd_sc_hd__a22o_1 _1749_ (.A1(_0557_),
    .A2(net182),
    .B1(_0445_),
    .B2(_0546_),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_4 _1750_ (.A(_0412_),
    .X(_0558_));
 sky130_fd_sc_hd__and3b_1 _1751_ (.A_N(_0451_),
    .B(_0558_),
    .C(net10),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _1752_ (.A1(_0450_),
    .A2(_0559_),
    .B1(_0557_),
    .B2(net103),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_1 _1753_ (.A1(_0557_),
    .A2(net200),
    .B1(_0519_),
    .B2(_0546_),
    .X(_0092_));
 sky130_fd_sc_hd__and3b_1 _1754_ (.A_N(_0451_),
    .B(_0558_),
    .C(net12),
    .X(_0560_));
 sky130_fd_sc_hd__a22o_1 _1755_ (.A1(_0450_),
    .A2(_0560_),
    .B1(_0557_),
    .B2(net120),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1756_ (.A0(_0427_),
    .A1(net339),
    .S(_0555_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_1 _1757_ (.A(_0561_),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _1758_ (.A1(_0557_),
    .A2(net202),
    .B1(_0453_),
    .B2(_0546_),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _1759_ (.A1(_0557_),
    .A2(net203),
    .B1(_0454_),
    .B2(_0546_),
    .X(_0096_));
 sky130_fd_sc_hd__nor2_1 _1760_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .B(_0543_),
    .Y(_0562_));
 sky130_fd_sc_hd__o2111ai_4 _1761_ (.A1(_0465_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0562_),
    .D1(_0928_),
    .Y(_0563_));
 sky130_fd_sc_hd__mux2_1 _1762_ (.A0(net8),
    .A1(net366),
    .S(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__clkbuf_1 _1763_ (.A(_0564_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _1764_ (.A0(_0419_),
    .A1(net270),
    .S(_0563_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1765_ (.A(_0565_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _1766_ (.A0(_0421_),
    .A1(net292),
    .S(_0563_),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_1 _1767_ (.A(_0566_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _1768_ (.A0(_0423_),
    .A1(net311),
    .S(_0563_),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _1769_ (.A(_0567_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _1770_ (.A0(_0425_),
    .A1(net305),
    .S(_0563_),
    .X(_0568_));
 sky130_fd_sc_hd__clkbuf_1 _1771_ (.A(_0568_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1772_ (.A0(_0427_),
    .A1(net343),
    .S(_0563_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_1 _1773_ (.A(_0569_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1774_ (.A0(_0429_),
    .A1(net322),
    .S(_0563_),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_1 _1775_ (.A(_0570_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1776_ (.A0(_0431_),
    .A1(net296),
    .S(_0563_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _1777_ (.A(_0571_),
    .X(_0104_));
 sky130_fd_sc_hd__o2111ai_4 _1778_ (.A1(_0465_),
    .A2(net35),
    .B1(_0410_),
    .C1(_0466_),
    .D1(_0545_),
    .Y(_0572_));
 sky130_fd_sc_hd__mux2_1 _1779_ (.A0(net8),
    .A1(net304),
    .S(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__clkbuf_1 _1780_ (.A(_0573_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1781_ (.A0(_0419_),
    .A1(net308),
    .S(_0572_),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_1 _1782_ (.A(_0574_),
    .X(_0106_));
 sky130_fd_sc_hd__a32o_1 _1783_ (.A1(_0473_),
    .A2(_0466_),
    .A3(_0559_),
    .B1(_0572_),
    .B2(net73),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(_0423_),
    .A1(net345),
    .S(_0572_),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_1 _1785_ (.A(_0575_),
    .X(_0108_));
 sky130_fd_sc_hd__a32o_1 _1786_ (.A1(_0473_),
    .A2(_0466_),
    .A3(_0560_),
    .B1(_0572_),
    .B2(net142),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1787_ (.A0(_0427_),
    .A1(net298),
    .S(_0572_),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_1 _1788_ (.A(_0576_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1789_ (.A0(_0429_),
    .A1(net293),
    .S(_0572_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _1790_ (.A(_0577_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1791_ (.A0(net15),
    .A1(net331),
    .S(_0572_),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_1 _1792_ (.A(_0578_),
    .X(_0112_));
 sky130_fd_sc_hd__buf_4 _1793_ (.A(_0523_),
    .X(_0579_));
 sky130_fd_sc_hd__nand4_2 _1794_ (.A(_0441_),
    .B(_0443_),
    .C(_0439_),
    .D(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__and4_1 _1795_ (.A(_0506_),
    .B(_0416_),
    .C(net8),
    .D(_0444_),
    .X(_0581_));
 sky130_fd_sc_hd__a22o_1 _1796_ (.A1(net198),
    .A2(_0580_),
    .B1(_0581_),
    .B2(_0579_),
    .X(_0113_));
 sky130_fd_sc_hd__o31a_1 _1797_ (.A1(_0451_),
    .A2(_0558_),
    .A3(_0503_),
    .B1(net321),
    .X(_0582_));
 sky130_fd_sc_hd__a31o_1 _1798_ (.A1(_0419_),
    .A2(_0502_),
    .A3(_0579_),
    .B1(_0582_),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_1 _1799_ (.A1(_0580_),
    .A2(net195),
    .B1(_0509_),
    .B2(_0579_),
    .X(_0115_));
 sky130_fd_sc_hd__and4_1 _1800_ (.A(_0506_),
    .B(_0416_),
    .C(net11),
    .D(_0444_),
    .X(_0583_));
 sky130_fd_sc_hd__a22o_1 _1801_ (.A1(net174),
    .A2(_0580_),
    .B1(_0583_),
    .B2(_0579_),
    .X(_0116_));
 sky130_fd_sc_hd__o31a_1 _1802_ (.A1(_0451_),
    .A2(_0558_),
    .A3(_0503_),
    .B1(net231),
    .X(_0584_));
 sky130_fd_sc_hd__a31o_1 _1803_ (.A1(_0425_),
    .A2(_0502_),
    .A3(_0579_),
    .B1(_0584_),
    .X(_0117_));
 sky130_fd_sc_hd__o31a_1 _1804_ (.A1(_0451_),
    .A2(_0558_),
    .A3(_0503_),
    .B1(net225),
    .X(_0585_));
 sky130_fd_sc_hd__a31o_1 _1805_ (.A1(_0427_),
    .A2(_0502_),
    .A3(_0579_),
    .B1(_0585_),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_1 _1806_ (.A1(_0580_),
    .A2(net230),
    .B1(_0513_),
    .B2(_0579_),
    .X(_0119_));
 sky130_fd_sc_hd__o31a_1 _1807_ (.A1(_0451_),
    .A2(_0558_),
    .A3(_0503_),
    .B1(net236),
    .X(_0586_));
 sky130_fd_sc_hd__a31o_1 _1808_ (.A1(_0431_),
    .A2(_0502_),
    .A3(_0579_),
    .B1(_0586_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_4 _1809_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[0] ),
    .X(_0587_));
 sky130_fd_sc_hd__o22ai_2 _1810_ (.A1(_0976_),
    .A2(_0977_),
    .B1(_0978_),
    .B2(_0979_),
    .Y(_0588_));
 sky130_fd_sc_hd__clkbuf_8 _1811_ (.A(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__o221ai_4 _1812_ (.A1(_0970_),
    .A2(_0971_),
    .B1(_0973_),
    .B2(_0974_),
    .C1(_0476_),
    .Y(_0590_));
 sky130_fd_sc_hd__and2_1 _1813_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[0] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tvalid_reg ),
    .X(_0591_));
 sky130_fd_sc_hd__clkbuf_4 _1814_ (.A(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__clkinv_4 _1815_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[2] ),
    .Y(_0593_));
 sky130_fd_sc_hd__nor2_2 _1816_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .B(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__o2111a_4 _1817_ (.A1(_0589_),
    .A2(net34),
    .B1(_0592_),
    .C1(_0594_),
    .D1(_0972_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _1818_ (.A0(net261),
    .A1(_0587_),
    .S(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_1 _1819_ (.A(_0596_),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_4 _1820_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[1] ),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _1821_ (.A0(net250),
    .A1(_0597_),
    .S(_0595_),
    .X(_0598_));
 sky130_fd_sc_hd__clkbuf_1 _1822_ (.A(_0598_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1823_ (.A0(net273),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ),
    .S(_0595_),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_1 _1824_ (.A(_0599_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1825_ (.A0(net255),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ),
    .S(_0595_),
    .X(_0600_));
 sky130_fd_sc_hd__clkbuf_1 _1826_ (.A(_0600_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_4 _1827_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[4] ),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _1828_ (.A0(net278),
    .A1(_0601_),
    .S(_0595_),
    .X(_0602_));
 sky130_fd_sc_hd__clkbuf_1 _1829_ (.A(_0602_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _1830_ (.A0(net252),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ),
    .S(_0595_),
    .X(_0603_));
 sky130_fd_sc_hd__clkbuf_1 _1831_ (.A(_0603_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(net266),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ),
    .S(_0595_),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_1 _1833_ (.A(_0604_),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_4 _1834_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[7] ),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _1835_ (.A0(net245),
    .A1(_0605_),
    .S(_0595_),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_1 _1836_ (.A(_0606_),
    .X(_0128_));
 sky130_fd_sc_hd__o2111ai_4 _1837_ (.A1(_0465_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0435_),
    .D1(_0523_),
    .Y(_0607_));
 sky130_fd_sc_hd__mux2_1 _1838_ (.A0(net8),
    .A1(net282),
    .S(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_1 _1839_ (.A(_0608_),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_1 _1840_ (.A1(_0607_),
    .A2(net199),
    .B1(_0445_),
    .B2(_0579_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1841_ (.A0(_0421_),
    .A1(net344),
    .S(_0607_),
    .X(_0609_));
 sky130_fd_sc_hd__clkbuf_1 _1842_ (.A(_0609_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1843_ (.A0(net11),
    .A1(net276),
    .S(_0607_),
    .X(_0610_));
 sky130_fd_sc_hd__clkbuf_1 _1844_ (.A(_0610_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1845_ (.A0(net12),
    .A1(net362),
    .S(_0607_),
    .X(_0611_));
 sky130_fd_sc_hd__clkbuf_1 _1846_ (.A(_0611_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1847_ (.A0(net13),
    .A1(net354),
    .S(_0607_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_1 _1848_ (.A(_0612_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1849_ (.A0(_0429_),
    .A1(net286),
    .S(_0607_),
    .X(_0613_));
 sky130_fd_sc_hd__clkbuf_1 _1850_ (.A(_0613_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _1851_ (.A0(net15),
    .A1(net361),
    .S(_0607_),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_1 _1852_ (.A(_0614_),
    .X(_0136_));
 sky130_fd_sc_hd__nor3_1 _1853_ (.A(_0413_),
    .B(_0412_),
    .C(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ),
    .Y(_0615_));
 sky130_fd_sc_hd__o2111ai_4 _1854_ (.A1(_0465_),
    .A2(_0407_),
    .B1(_0411_),
    .C1(_0615_),
    .D1(_0928_),
    .Y(_0616_));
 sky130_fd_sc_hd__mux2_1 _1855_ (.A0(net8),
    .A1(net330),
    .S(net28),
    .X(_0617_));
 sky130_fd_sc_hd__clkbuf_1 _1856_ (.A(_0617_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1857_ (.A0(net9),
    .A1(net347),
    .S(net28),
    .X(_0618_));
 sky130_fd_sc_hd__clkbuf_1 _1858_ (.A(_0618_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _1859_ (.A0(net10),
    .A1(net358),
    .S(net28),
    .X(_0619_));
 sky130_fd_sc_hd__clkbuf_1 _1860_ (.A(_0619_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _1861_ (.A0(net11),
    .A1(net303),
    .S(net28),
    .X(_0620_));
 sky130_fd_sc_hd__clkbuf_1 _1862_ (.A(_0620_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _1863_ (.A0(net12),
    .A1(net365),
    .S(_0616_),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_1 _1864_ (.A(_0621_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _1865_ (.A0(net13),
    .A1(net364),
    .S(_0616_),
    .X(_0622_));
 sky130_fd_sc_hd__clkbuf_1 _1866_ (.A(_0622_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _1867_ (.A0(net14),
    .A1(net359),
    .S(_0616_),
    .X(_0623_));
 sky130_fd_sc_hd__clkbuf_1 _1868_ (.A(_0623_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _1869_ (.A0(net15),
    .A1(net368),
    .S(_0616_),
    .X(_0624_));
 sky130_fd_sc_hd__clkbuf_1 _1870_ (.A(_0624_),
    .X(_0144_));
 sky130_fd_sc_hd__nand2_4 _1871_ (.A(_0434_),
    .B(_0501_),
    .Y(_0625_));
 sky130_fd_sc_hd__a22o_1 _1872_ (.A1(net194),
    .A2(_0625_),
    .B1(_0581_),
    .B2(_0446_),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_1 _1873_ (.A1(net132),
    .A2(_0625_),
    .B1(_0508_),
    .B2(_0446_),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _1874_ (.A1(net172),
    .A2(_0625_),
    .B1(_0509_),
    .B2(_0446_),
    .X(_0147_));
 sky130_fd_sc_hd__a22o_1 _1875_ (.A1(net155),
    .A2(_0625_),
    .B1(_0583_),
    .B2(_0446_),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_1 _1876_ (.A1(net210),
    .A2(_0625_),
    .B1(_0511_),
    .B2(_0446_),
    .X(_0149_));
 sky130_fd_sc_hd__a22o_1 _1877_ (.A1(net143),
    .A2(_0625_),
    .B1(_0512_),
    .B2(_0446_),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _1878_ (.A1(net164),
    .A2(_0625_),
    .B1(_0513_),
    .B2(_0446_),
    .X(_0151_));
 sky130_fd_sc_hd__a31o_1 _1879_ (.A1(_0451_),
    .A2(_0558_),
    .A3(_0501_),
    .B1(net240),
    .X(_0626_));
 sky130_fd_sc_hd__o21a_1 _1880_ (.A1(_0431_),
    .A2(_0625_),
    .B1(_0626_),
    .X(_0152_));
 sky130_fd_sc_hd__and2_2 _1881_ (.A(_0593_),
    .B(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .X(_0627_));
 sky130_fd_sc_hd__inv_2 _1882_ (.A(_0972_),
    .Y(_0628_));
 sky130_fd_sc_hd__o2111a_4 _1883_ (.A1(_0589_),
    .A2(_0590_),
    .B1(_0592_),
    .C1(_0627_),
    .D1(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _1884_ (.A0(net246),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[0] ),
    .S(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__clkbuf_1 _1885_ (.A(_0630_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _1886_ (.A0(net251),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[1] ),
    .S(_0629_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _1887_ (.A(_0631_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _1888_ (.A0(net244),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ),
    .S(_0629_),
    .X(_0632_));
 sky130_fd_sc_hd__clkbuf_1 _1889_ (.A(_0632_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _1890_ (.A0(net288),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ),
    .S(_0629_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _1891_ (.A(_0633_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _1892_ (.A0(net259),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[4] ),
    .S(_0629_),
    .X(_0634_));
 sky130_fd_sc_hd__clkbuf_1 _1893_ (.A(_0634_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1894_ (.A0(net256),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ),
    .S(_0629_),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_1 _1895_ (.A(_0635_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _1896_ (.A0(net249),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ),
    .S(_0629_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_1 _1897_ (.A(_0636_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _1898_ (.A0(net262),
    .A1(_0605_),
    .S(_0629_),
    .X(_0637_));
 sky130_fd_sc_hd__clkbuf_1 _1899_ (.A(_0637_),
    .X(_0160_));
 sky130_fd_sc_hd__buf_4 _1900_ (.A(_0594_),
    .X(_0638_));
 sky130_fd_sc_hd__inv_2 _1901_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[0] ),
    .Y(_0639_));
 sky130_fd_sc_hd__o2111a_1 _1902_ (.A1(_0589_),
    .A2(_0590_),
    .B1(_0972_),
    .C1(_0639_),
    .D1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tvalid_reg ),
    .X(_0640_));
 sky130_fd_sc_hd__buf_4 _1903_ (.A(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__buf_4 _1904_ (.A(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__buf_4 _1905_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .X(_0643_));
 sky130_fd_sc_hd__nand3b_4 _1906_ (.A_N(_0643_),
    .B(_0479_),
    .C(_0641_),
    .Y(_0644_));
 sky130_fd_sc_hd__a32o_1 _1907_ (.A1(_0587_),
    .A2(_0638_),
    .A3(_0642_),
    .B1(_0644_),
    .B2(net167),
    .X(_0161_));
 sky130_fd_sc_hd__a32o_1 _1908_ (.A1(_0597_),
    .A2(_0638_),
    .A3(_0642_),
    .B1(_0644_),
    .B2(net168),
    .X(_0162_));
 sky130_fd_sc_hd__a32o_1 _1909_ (.A1(_0489_),
    .A2(_0638_),
    .A3(_0642_),
    .B1(_0644_),
    .B2(net71),
    .X(_0163_));
 sky130_fd_sc_hd__a32o_1 _1910_ (.A1(_0491_),
    .A2(_0638_),
    .A3(_0642_),
    .B1(_0644_),
    .B2(net84),
    .X(_0164_));
 sky130_fd_sc_hd__a32o_1 _1911_ (.A1(_0601_),
    .A2(_0638_),
    .A3(_0642_),
    .B1(_0644_),
    .B2(net74),
    .X(_0165_));
 sky130_fd_sc_hd__a32o_1 _1912_ (.A1(_0494_),
    .A2(_0638_),
    .A3(_0642_),
    .B1(_0644_),
    .B2(net105),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_4 _1913_ (.A(_0594_),
    .X(_0645_));
 sky130_fd_sc_hd__a32o_1 _1914_ (.A1(_0496_),
    .A2(_0645_),
    .A3(_0642_),
    .B1(_0644_),
    .B2(net89),
    .X(_0167_));
 sky130_fd_sc_hd__a32o_1 _1915_ (.A1(_0605_),
    .A2(_0645_),
    .A3(_0642_),
    .B1(_0644_),
    .B2(net69),
    .X(_0168_));
 sky130_fd_sc_hd__buf_4 _1916_ (.A(_0628_),
    .X(_0646_));
 sky130_fd_sc_hd__nand3_4 _1917_ (.A(_0476_),
    .B(_0975_),
    .C(_0980_),
    .Y(_0647_));
 sky130_fd_sc_hd__buf_4 _1918_ (.A(_0592_),
    .X(_0648_));
 sky130_fd_sc_hd__nand4_4 _1919_ (.A(_0646_),
    .B(_0647_),
    .C(_0648_),
    .D(_0594_),
    .Y(_0649_));
 sky130_fd_sc_hd__and3_1 _1920_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[0] ),
    .B(_0483_),
    .C(_0646_),
    .X(_0650_));
 sky130_fd_sc_hd__a22o_1 _1921_ (.A1(net156),
    .A2(_0649_),
    .B1(_0650_),
    .B2(_0638_),
    .X(_0169_));
 sky130_fd_sc_hd__and3_1 _1922_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[1] ),
    .B(_0483_),
    .C(_0646_),
    .X(_0651_));
 sky130_fd_sc_hd__a22o_1 _1923_ (.A1(net162),
    .A2(_0649_),
    .B1(_0651_),
    .B2(_0638_),
    .X(_0170_));
 sky130_fd_sc_hd__or2_2 _1924_ (.A(_0643_),
    .B(_0593_),
    .X(_0652_));
 sky130_fd_sc_hd__o2111ai_2 _1925_ (.A1(_0589_),
    .A2(net34),
    .B1(_0648_),
    .C1(_0646_),
    .D1(_0489_),
    .Y(_0653_));
 sky130_fd_sc_hd__a2bb2o_1 _1926_ (.A1_N(_0652_),
    .A2_N(_0653_),
    .B1(_0649_),
    .B2(net184),
    .X(_0171_));
 sky130_fd_sc_hd__o2111ai_4 _1927_ (.A1(_0589_),
    .A2(net34),
    .B1(_0648_),
    .C1(_0646_),
    .D1(_0491_),
    .Y(_0654_));
 sky130_fd_sc_hd__a2bb2o_1 _1928_ (.A1_N(_0652_),
    .A2_N(_0654_),
    .B1(_0649_),
    .B2(net117),
    .X(_0172_));
 sky130_fd_sc_hd__and3_1 _1929_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[4] ),
    .B(_0478_),
    .C(_0646_),
    .X(_0655_));
 sky130_fd_sc_hd__a22o_1 _1930_ (.A1(net136),
    .A2(_0649_),
    .B1(_0655_),
    .B2(_0638_),
    .X(_0173_));
 sky130_fd_sc_hd__o2111ai_2 _1931_ (.A1(_0589_),
    .A2(net34),
    .B1(_0648_),
    .C1(_0646_),
    .D1(_0494_),
    .Y(_0656_));
 sky130_fd_sc_hd__a2bb2o_1 _1932_ (.A1_N(_0652_),
    .A2_N(_0656_),
    .B1(_0649_),
    .B2(net126),
    .X(_0174_));
 sky130_fd_sc_hd__o2111ai_2 _1933_ (.A1(_0589_),
    .A2(net34),
    .B1(_0648_),
    .C1(_0646_),
    .D1(_0496_),
    .Y(_0657_));
 sky130_fd_sc_hd__a2bb2o_1 _1934_ (.A1_N(_0652_),
    .A2_N(_0657_),
    .B1(_0649_),
    .B2(net116),
    .X(_0175_));
 sky130_fd_sc_hd__and3_1 _1935_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[7] ),
    .B(_0478_),
    .C(_0646_),
    .X(_0658_));
 sky130_fd_sc_hd__a22o_1 _1936_ (.A1(net144),
    .A2(_0649_),
    .B1(_0658_),
    .B2(_0638_),
    .X(_0176_));
 sky130_fd_sc_hd__o2111a_1 _1937_ (.A1(_0588_),
    .A2(_0590_),
    .B1(_0628_),
    .C1(_0639_),
    .D1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tvalid_reg ),
    .X(_0659_));
 sky130_fd_sc_hd__buf_4 _1938_ (.A(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__buf_4 _1939_ (.A(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__nand3b_4 _1940_ (.A_N(_0643_),
    .B(_0479_),
    .C(_0660_),
    .Y(_0662_));
 sky130_fd_sc_hd__a32o_1 _1941_ (.A1(_0587_),
    .A2(_0645_),
    .A3(_0661_),
    .B1(_0662_),
    .B2(net110),
    .X(_0177_));
 sky130_fd_sc_hd__a32o_1 _1942_ (.A1(_0597_),
    .A2(_0645_),
    .A3(_0661_),
    .B1(_0662_),
    .B2(net77),
    .X(_0178_));
 sky130_fd_sc_hd__a32o_1 _1943_ (.A1(_0489_),
    .A2(_0645_),
    .A3(_0661_),
    .B1(_0662_),
    .B2(net137),
    .X(_0179_));
 sky130_fd_sc_hd__a32o_1 _1944_ (.A1(_0491_),
    .A2(_0645_),
    .A3(_0661_),
    .B1(_0662_),
    .B2(net86),
    .X(_0180_));
 sky130_fd_sc_hd__a32o_1 _1945_ (.A1(_0601_),
    .A2(_0645_),
    .A3(_0661_),
    .B1(_0662_),
    .B2(net87),
    .X(_0181_));
 sky130_fd_sc_hd__a32o_1 _1946_ (.A1(_0494_),
    .A2(_0645_),
    .A3(_0661_),
    .B1(_0662_),
    .B2(net76),
    .X(_0182_));
 sky130_fd_sc_hd__a32o_1 _1947_ (.A1(_0496_),
    .A2(_0645_),
    .A3(_0661_),
    .B1(_0662_),
    .B2(net88),
    .X(_0183_));
 sky130_fd_sc_hd__a32o_1 _1948_ (.A1(_0605_),
    .A2(_0645_),
    .A3(_0661_),
    .B1(_0662_),
    .B2(net68),
    .X(_0184_));
 sky130_fd_sc_hd__and3_1 _1949_ (.A(_0647_),
    .B(_0592_),
    .C(_0972_),
    .X(_0663_));
 sky130_fd_sc_hd__nor2_2 _1950_ (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .B(_0479_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_4 _1951_ (.A(_0663_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__clkbuf_4 _1952_ (.A(_0664_),
    .X(_0666_));
 sky130_fd_sc_hd__clkbuf_4 _1953_ (.A(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__a22o_1 _1954_ (.A1(_0665_),
    .A2(net177),
    .B1(_0484_),
    .B2(_0667_),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _1955_ (.A1(_0665_),
    .A2(net201),
    .B1(_0488_),
    .B2(_0667_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _1956_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ),
    .B(_0482_),
    .C(_0483_),
    .X(_0668_));
 sky130_fd_sc_hd__a22o_1 _1957_ (.A1(_0667_),
    .A2(_0668_),
    .B1(_0665_),
    .B2(net178),
    .X(_0187_));
 sky130_fd_sc_hd__and3_1 _1958_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ),
    .B(_0482_),
    .C(_0483_),
    .X(_0669_));
 sky130_fd_sc_hd__a22o_1 _1959_ (.A1(_0667_),
    .A2(_0669_),
    .B1(_0665_),
    .B2(net165),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_1 _1960_ (.A1(_0665_),
    .A2(net179),
    .B1(_0493_),
    .B2(_0667_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_4 _1961_ (.A(_0666_),
    .X(_0670_));
 sky130_fd_sc_hd__and3_1 _1962_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ),
    .B(_0482_),
    .C(_0483_),
    .X(_0671_));
 sky130_fd_sc_hd__a22o_1 _1963_ (.A1(_0670_),
    .A2(_0671_),
    .B1(_0665_),
    .B2(net134),
    .X(_0190_));
 sky130_fd_sc_hd__and3_1 _1964_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ),
    .B(_0482_),
    .C(_0483_),
    .X(_0672_));
 sky130_fd_sc_hd__a22o_1 _1965_ (.A1(_0670_),
    .A2(_0672_),
    .B1(_0665_),
    .B2(net140),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _1966_ (.A1(_0665_),
    .A2(net181),
    .B1(_0498_),
    .B2(_0667_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_4 _1967_ (.A(_0641_),
    .X(_0673_));
 sky130_fd_sc_hd__nand3b_4 _1968_ (.A_N(_0643_),
    .B(_0641_),
    .C(_0593_),
    .Y(_0674_));
 sky130_fd_sc_hd__a32o_1 _1969_ (.A1(_0587_),
    .A2(_0673_),
    .A3(_0670_),
    .B1(_0674_),
    .B2(net118),
    .X(_0193_));
 sky130_fd_sc_hd__a32o_1 _1970_ (.A1(_0597_),
    .A2(_0673_),
    .A3(_0670_),
    .B1(_0674_),
    .B2(net125),
    .X(_0194_));
 sky130_fd_sc_hd__a32o_1 _1971_ (.A1(_0489_),
    .A2(_0673_),
    .A3(_0670_),
    .B1(_0674_),
    .B2(net98),
    .X(_0195_));
 sky130_fd_sc_hd__a32o_1 _1972_ (.A1(_0491_),
    .A2(_0673_),
    .A3(_0670_),
    .B1(_0674_),
    .B2(net82),
    .X(_0196_));
 sky130_fd_sc_hd__a32o_1 _1973_ (.A1(_0601_),
    .A2(_0673_),
    .A3(_0670_),
    .B1(_0674_),
    .B2(net75),
    .X(_0197_));
 sky130_fd_sc_hd__a32o_1 _1974_ (.A1(_0494_),
    .A2(_0673_),
    .A3(_0670_),
    .B1(_0674_),
    .B2(net130),
    .X(_0198_));
 sky130_fd_sc_hd__a32o_1 _1975_ (.A1(_0496_),
    .A2(_0641_),
    .A3(_0670_),
    .B1(_0674_),
    .B2(net119),
    .X(_0199_));
 sky130_fd_sc_hd__a32o_1 _1976_ (.A1(_0605_),
    .A2(_0641_),
    .A3(_0670_),
    .B1(_0674_),
    .B2(net113),
    .X(_0200_));
 sky130_fd_sc_hd__nand4_4 _1977_ (.A(_0646_),
    .B(_0647_),
    .C(_0648_),
    .D(_0664_),
    .Y(_0675_));
 sky130_fd_sc_hd__a22o_1 _1978_ (.A1(_0675_),
    .A2(net185),
    .B1(_0650_),
    .B2(_0667_),
    .X(_0201_));
 sky130_fd_sc_hd__a22o_1 _1979_ (.A1(_0675_),
    .A2(net183),
    .B1(_0651_),
    .B2(_0667_),
    .X(_0202_));
 sky130_fd_sc_hd__or2_1 _1980_ (.A(_0643_),
    .B(_0479_),
    .X(_0676_));
 sky130_fd_sc_hd__a2bb2o_1 _1981_ (.A1_N(_0653_),
    .A2_N(_0676_),
    .B1(_0675_),
    .B2(net147),
    .X(_0203_));
 sky130_fd_sc_hd__a2bb2o_1 _1982_ (.A1_N(_0654_),
    .A2_N(_0676_),
    .B1(_0675_),
    .B2(net135),
    .X(_0204_));
 sky130_fd_sc_hd__a22o_1 _1983_ (.A1(_0675_),
    .A2(net191),
    .B1(_0655_),
    .B2(_0667_),
    .X(_0205_));
 sky130_fd_sc_hd__a2bb2o_1 _1984_ (.A1_N(_0656_),
    .A2_N(_0676_),
    .B1(_0675_),
    .B2(net131),
    .X(_0206_));
 sky130_fd_sc_hd__a2bb2o_1 _1985_ (.A1_N(_0657_),
    .A2_N(_0676_),
    .B1(_0675_),
    .B2(net129),
    .X(_0207_));
 sky130_fd_sc_hd__a22o_1 _1986_ (.A1(_0675_),
    .A2(net190),
    .B1(_0658_),
    .B2(_0667_),
    .X(_0208_));
 sky130_fd_sc_hd__clkinv_4 _1987_ (.A(net6),
    .Y(_0677_));
 sky130_fd_sc_hd__clkbuf_4 _1988_ (.A(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__and4b_2 _1989_ (.A_N(net16),
    .B(net5),
    .C(net7),
    .D(net41),
    .X(_0679_));
 sky130_fd_sc_hd__a21oi_1 _1990_ (.A1(_0981_),
    .A2(_0679_),
    .B1(_0986_),
    .Y(_0680_));
 sky130_fd_sc_hd__o22ai_1 _1991_ (.A1(_0970_),
    .A2(_0971_),
    .B1(_0973_),
    .B2(_0974_),
    .Y(_0681_));
 sky130_fd_sc_hd__o311a_1 _1992_ (.A1(_0476_),
    .A2(_0681_),
    .A3(_0589_),
    .B1(_0679_),
    .C1(_0986_),
    .X(_0682_));
 sky130_fd_sc_hd__nor3_1 _1993_ (.A(_0678_),
    .B(_0680_),
    .C(_0682_),
    .Y(_0209_));
 sky130_fd_sc_hd__a31o_1 _1994_ (.A1(_0981_),
    .A2(_0679_),
    .A3(_0986_),
    .B1(_0987_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_4 _1995_ (.A(_1037_),
    .X(_0684_));
 sky130_fd_sc_hd__nand4_2 _1996_ (.A(_0981_),
    .B(_0679_),
    .C(_0987_),
    .D(_0986_),
    .Y(_0685_));
 sky130_fd_sc_hd__and3_1 _1997_ (.A(_0683_),
    .B(_0684_),
    .C(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_1 _1998_ (.A(_0686_),
    .X(_0210_));
 sky130_fd_sc_hd__a31o_1 _1999_ (.A1(_0947_),
    .A2(_0987_),
    .A3(_0682_),
    .B1(_0677_),
    .X(_0687_));
 sky130_fd_sc_hd__a21oi_1 _2000_ (.A1(_0960_),
    .A2(_0685_),
    .B1(_0687_),
    .Y(_0211_));
 sky130_fd_sc_hd__and2_1 _2001_ (.A(_0947_),
    .B(_0987_),
    .X(_0688_));
 sky130_fd_sc_hd__buf_4 _2002_ (.A(_0677_),
    .X(_0689_));
 sky130_fd_sc_hd__o21a_1 _2003_ (.A1(_0960_),
    .A2(_0685_),
    .B1(_0942_),
    .X(_0690_));
 sky130_fd_sc_hd__a311oi_1 _2004_ (.A1(_0951_),
    .A2(_0682_),
    .A3(_0688_),
    .B1(_0689_),
    .C1(_0690_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor3_1 _2005_ (.A(_0942_),
    .B(_0960_),
    .C(_0685_),
    .Y(_0691_));
 sky130_fd_sc_hd__nand4_1 _2006_ (.A(net357),
    .B(_0951_),
    .C(_0682_),
    .D(_0688_),
    .Y(_0692_));
 sky130_fd_sc_hd__clkbuf_4 _2007_ (.A(_0684_),
    .X(_0693_));
 sky130_fd_sc_hd__o211a_1 _2008_ (.A1(net357),
    .A2(_0691_),
    .B1(_0692_),
    .C1(_0693_),
    .X(_0213_));
 sky130_fd_sc_hd__a21oi_1 _2009_ (.A1(_0647_),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tvalid_reg ),
    .B1(net374),
    .Y(_0694_));
 sky130_fd_sc_hd__a211oi_1 _2010_ (.A1(_0647_),
    .A2(_0648_),
    .B1(_0689_),
    .C1(_0694_),
    .Y(_0214_));
 sky130_fd_sc_hd__a31o_1 _2011_ (.A1(_0647_),
    .A2(_0648_),
    .A3(_0482_),
    .B1(_0689_),
    .X(_0695_));
 sky130_fd_sc_hd__o21ba_1 _2012_ (.A1(_0482_),
    .A2(_0483_),
    .B1_N(_0695_),
    .X(_0215_));
 sky130_fd_sc_hd__a41o_1 _2013_ (.A1(_0647_),
    .A2(_0648_),
    .A3(_0479_),
    .A4(_0482_),
    .B1(_0677_),
    .X(_0696_));
 sky130_fd_sc_hd__o21ba_1 _2014_ (.A1(_0479_),
    .A2(_0663_),
    .B1_N(_0696_),
    .X(_0216_));
 sky130_fd_sc_hd__a31o_1 _2015_ (.A1(_0479_),
    .A2(_0972_),
    .A3(_0478_),
    .B1(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ),
    .X(_0697_));
 sky130_fd_sc_hd__and3_1 _2016_ (.A(_0697_),
    .B(_0684_),
    .C(_0481_),
    .X(_0698_));
 sky130_fd_sc_hd__clkbuf_1 _2017_ (.A(_0698_),
    .X(_0217_));
 sky130_fd_sc_hd__a31o_1 _2018_ (.A1(_0647_),
    .A2(_0592_),
    .A3(_0480_),
    .B1(\uart_inst.fifo_rx_inst.write_ptr_reg[4] ),
    .X(_0699_));
 sky130_fd_sc_hd__nand4_1 _2019_ (.A(_0647_),
    .B(_0648_),
    .C(_0480_),
    .D(\uart_inst.fifo_rx_inst.write_ptr_reg[4] ),
    .Y(_0700_));
 sky130_fd_sc_hd__and3_1 _2020_ (.A(_0699_),
    .B(_0684_),
    .C(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__clkbuf_1 _2021_ (.A(_0701_),
    .X(_0218_));
 sky130_fd_sc_hd__a41o_1 _2022_ (.A1(_1029_),
    .A2(_0939_),
    .A3(_0931_),
    .A4(_1034_),
    .B1(_0400_),
    .X(_0702_));
 sky130_fd_sc_hd__or3_1 _2023_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[3] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[2] ),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[1] ),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_1 _2024_ (.A(_0703_),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[0] ),
    .Y(_0704_));
 sky130_fd_sc_hd__a21oi_1 _2025_ (.A1(_1036_),
    .A2(_0704_),
    .B1(_0400_),
    .Y(_0705_));
 sky130_fd_sc_hd__a211o_1 _2026_ (.A1(_0702_),
    .A2(net356),
    .B1(_0678_),
    .C1(_0705_),
    .X(_0219_));
 sky130_fd_sc_hd__nor3_1 _2027_ (.A(_0934_),
    .B(_0401_),
    .C(_0465_),
    .Y(_0706_));
 sky130_fd_sc_hd__or3b_1 _2028_ (.A(_0706_),
    .B(_1075_),
    .C_N(\uart_inst.uart_core_inst.uart_tx_inst.s_axis_tready_reg ),
    .X(_0707_));
 sky130_fd_sc_hd__o2111a_1 _2029_ (.A1(net310),
    .A2(_1050_),
    .B1(_1091_),
    .C1(_0684_),
    .D1(_0707_),
    .X(_0220_));
 sky130_fd_sc_hd__nand3_4 _2030_ (.A(_0643_),
    .B(_0479_),
    .C(_0641_),
    .Y(_0708_));
 sky130_fd_sc_hd__a32o_1 _2031_ (.A1(_0587_),
    .A2(_0487_),
    .A3(_0642_),
    .B1(_0708_),
    .B2(net115),
    .X(_0221_));
 sky130_fd_sc_hd__a32o_1 _2032_ (.A1(_0597_),
    .A2(_0487_),
    .A3(_0642_),
    .B1(_0708_),
    .B2(net121),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_4 _2033_ (.A(_0641_),
    .X(_0709_));
 sky130_fd_sc_hd__a32o_1 _2034_ (.A1(_0489_),
    .A2(_0487_),
    .A3(_0709_),
    .B1(_0708_),
    .B2(net70),
    .X(_0223_));
 sky130_fd_sc_hd__a32o_1 _2035_ (.A1(_0491_),
    .A2(_0487_),
    .A3(_0709_),
    .B1(_0708_),
    .B2(net78),
    .X(_0224_));
 sky130_fd_sc_hd__buf_2 _2036_ (.A(_0486_),
    .X(_0710_));
 sky130_fd_sc_hd__a32o_1 _2037_ (.A1(_0601_),
    .A2(_0710_),
    .A3(_0709_),
    .B1(_0708_),
    .B2(net133),
    .X(_0225_));
 sky130_fd_sc_hd__a32o_1 _2038_ (.A1(_0494_),
    .A2(_0710_),
    .A3(_0709_),
    .B1(_0708_),
    .B2(net123),
    .X(_0226_));
 sky130_fd_sc_hd__a32o_1 _2039_ (.A1(_0496_),
    .A2(_0710_),
    .A3(_0709_),
    .B1(_0708_),
    .B2(net145),
    .X(_0227_));
 sky130_fd_sc_hd__a32o_1 _2040_ (.A1(_0605_),
    .A2(_0710_),
    .A3(_0709_),
    .B1(_0708_),
    .B2(net100),
    .X(_0228_));
 sky130_fd_sc_hd__o2111ai_4 _2041_ (.A1(_0589_),
    .A2(net34),
    .B1(_0592_),
    .C1(_0486_),
    .D1(_0628_),
    .Y(_0711_));
 sky130_fd_sc_hd__mux2_1 _2042_ (.A0(_0587_),
    .A1(net285),
    .S(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_1 _2043_ (.A(_0712_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2044_ (.A0(_0597_),
    .A1(net260),
    .S(_0711_),
    .X(_0713_));
 sky130_fd_sc_hd__clkbuf_1 _2045_ (.A(_0713_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2046_ (.A0(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ),
    .A1(net242),
    .S(_0711_),
    .X(_0714_));
 sky130_fd_sc_hd__clkbuf_1 _2047_ (.A(_0714_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2048_ (.A0(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ),
    .A1(net280),
    .S(_0711_),
    .X(_0715_));
 sky130_fd_sc_hd__clkbuf_1 _2049_ (.A(_0715_),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _2050_ (.A1(net187),
    .A2(_0711_),
    .B1(_0655_),
    .B2(_0487_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2051_ (.A0(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ),
    .A1(net327),
    .S(_0711_),
    .X(_0716_));
 sky130_fd_sc_hd__clkbuf_1 _2052_ (.A(_0716_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2053_ (.A0(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ),
    .A1(net268),
    .S(_0711_),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_1 _2054_ (.A(_0717_),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _2055_ (.A1(net141),
    .A2(_0711_),
    .B1(_0658_),
    .B2(_0487_),
    .X(_0236_));
 sky130_fd_sc_hd__o31a_1 _2056_ (.A1(_1042_),
    .A2(_1094_),
    .A3(_1041_),
    .B1(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[0] ),
    .X(_0718_));
 sky130_fd_sc_hd__o221ai_4 _2057_ (.A1(_0935_),
    .A2(_0936_),
    .B1(_0937_),
    .B2(_0938_),
    .C1(_1029_),
    .Y(_0719_));
 sky130_fd_sc_hd__o311a_1 _2058_ (.A1(_0403_),
    .A2(_0719_),
    .A3(_0703_),
    .B1(_1047_),
    .C1(_1032_),
    .X(_0720_));
 sky130_fd_sc_hd__o21a_1 _2059_ (.A1(_0718_),
    .A2(_0720_),
    .B1(_0693_),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_4 _2060_ (.A(_1037_),
    .X(_0721_));
 sky130_fd_sc_hd__nand4_1 _2061_ (.A(_1091_),
    .B(_1035_),
    .C(_1031_),
    .D(_1032_),
    .Y(_0722_));
 sky130_fd_sc_hd__o21ai_1 _2062_ (.A1(_1031_),
    .A2(_0720_),
    .B1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__o311a_1 _2063_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[3] ),
    .A2(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[2] ),
    .A3(net333),
    .B1(_0721_),
    .C1(_0723_),
    .X(_0238_));
 sky130_fd_sc_hd__a41o_1 _2064_ (.A1(_1091_),
    .A2(_1035_),
    .A3(_1031_),
    .A4(_1032_),
    .B1(_1030_),
    .X(_0724_));
 sky130_fd_sc_hd__o311a_1 _2065_ (.A1(_0403_),
    .A2(_0719_),
    .A3(_0703_),
    .B1(_1047_),
    .C1(_1032_),
    .X(_0725_));
 sky130_fd_sc_hd__nand4_1 _2066_ (.A(_1030_),
    .B(_0725_),
    .C(_1031_),
    .D(net351),
    .Y(_0726_));
 sky130_fd_sc_hd__a21oi_1 _2067_ (.A1(_0724_),
    .A2(_0726_),
    .B1(_0678_),
    .Y(_0239_));
 sky130_fd_sc_hd__a311o_1 _2068_ (.A1(_1029_),
    .A2(_0939_),
    .A3(_0931_),
    .B1(_0400_),
    .C1(_1075_),
    .X(_0727_));
 sky130_fd_sc_hd__o21ai_1 _2069_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[2] ),
    .A2(_0722_),
    .B1(net351),
    .Y(_0728_));
 sky130_fd_sc_hd__a21oi_1 _2070_ (.A1(_0727_),
    .A2(_0728_),
    .B1(_0678_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand3_2 _2071_ (.A(_1047_),
    .B(net27),
    .C(_1034_),
    .Y(_0729_));
 sky130_fd_sc_hd__a21oi_1 _2072_ (.A1(_1097_),
    .A2(_0729_),
    .B1(net337),
    .Y(_0730_));
 sky130_fd_sc_hd__a31o_1 _2073_ (.A1(_1097_),
    .A2(_0729_),
    .A3(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ),
    .B1(_0677_),
    .X(_0731_));
 sky130_fd_sc_hd__nor2_1 _2074_ (.A(_0730_),
    .B(_0731_),
    .Y(_0242_));
 sky130_fd_sc_hd__or3_1 _2075_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[2] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[0] ),
    .X(_0732_));
 sky130_fd_sc_hd__o21ai_1 _2076_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ),
    .A2(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[0] ),
    .B1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[2] ),
    .Y(_0733_));
 sky130_fd_sc_hd__a21o_1 _2077_ (.A1(_0732_),
    .A2(_0733_),
    .B1(_1091_),
    .X(_0734_));
 sky130_fd_sc_hd__nor2_1 _2078_ (.A(_0400_),
    .B(_1035_),
    .Y(_0735_));
 sky130_fd_sc_hd__a211oi_1 _2079_ (.A1(_1096_),
    .A2(_0734_),
    .B1(_0735_),
    .C1(_0689_),
    .Y(_0243_));
 sky130_fd_sc_hd__o31a_1 _2080_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[2] ),
    .A2(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ),
    .A3(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[0] ),
    .B1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[3] ),
    .X(_0736_));
 sky130_fd_sc_hd__o21ai_1 _2081_ (.A1(net39),
    .A2(_0736_),
    .B1(_0400_),
    .Y(_0737_));
 sky130_fd_sc_hd__a211oi_1 _2082_ (.A1(_1096_),
    .A2(_0737_),
    .B1(_0689_),
    .C1(_0735_),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _2083_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[4] ),
    .Y(_0738_));
 sky130_fd_sc_hd__xor2_1 _2084_ (.A(_0738_),
    .B(net39),
    .X(_0739_));
 sky130_fd_sc_hd__o21ai_1 _2085_ (.A1(_1091_),
    .A2(_0739_),
    .B1(_1096_),
    .Y(_0740_));
 sky130_fd_sc_hd__o311a_1 _2086_ (.A1(_0400_),
    .A2(_1090_),
    .A3(_1075_),
    .B1(_0721_),
    .C1(_0740_),
    .X(_0245_));
 sky130_fd_sc_hd__or4_1 _2087_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[3] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[2] ),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ),
    .D(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[0] ),
    .X(_0741_));
 sky130_fd_sc_hd__or3_1 _2088_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[5] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[4] ),
    .C(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__o21ai_1 _2089_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[4] ),
    .A2(_0741_),
    .B1(net332),
    .Y(_0743_));
 sky130_fd_sc_hd__a221oi_1 _2090_ (.A1(_1036_),
    .A2(_1091_),
    .B1(_0742_),
    .B2(_0743_),
    .C1(_0689_),
    .Y(_0246_));
 sky130_fd_sc_hd__nor2_1 _2091_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[5] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[4] ),
    .Y(_0744_));
 sky130_fd_sc_hd__a31oi_1 _2092_ (.A1(_0729_),
    .A2(_0744_),
    .A3(net376),
    .B1(net217),
    .Y(_0745_));
 sky130_fd_sc_hd__a311oi_1 _2093_ (.A1(net217),
    .A2(net376),
    .A3(_0744_),
    .B1(_0689_),
    .C1(_0745_),
    .Y(_0247_));
 sky130_fd_sc_hd__buf_2 _2094_ (.A(_0399_),
    .X(_0746_));
 sky130_fd_sc_hd__o41ai_1 _2095_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[6] ),
    .A2(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[5] ),
    .A3(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[4] ),
    .A4(_0741_),
    .B1(net204),
    .Y(_0747_));
 sky130_fd_sc_hd__a41o_2 _2096_ (.A1(net39),
    .A2(net375),
    .A3(_1095_),
    .A4(_1040_),
    .B1(_0677_),
    .X(_0748_));
 sky130_fd_sc_hd__a21oi_1 _2097_ (.A1(_0746_),
    .A2(net205),
    .B1(_0748_),
    .Y(_0248_));
 sky130_fd_sc_hd__o21ai_1 _2098_ (.A1(_0746_),
    .A2(_0735_),
    .B1(net371),
    .Y(_0749_));
 sky130_fd_sc_hd__a311o_1 _2099_ (.A1(_1091_),
    .A2(net27),
    .A3(_1034_),
    .B1(_0746_),
    .C1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[8] ),
    .X(_0750_));
 sky130_fd_sc_hd__a21oi_1 _2100_ (.A1(_0749_),
    .A2(_0750_),
    .B1(_0678_),
    .Y(_0249_));
 sky130_fd_sc_hd__o21bai_1 _2101_ (.A1(_0400_),
    .A2(_1035_),
    .B1_N(_0746_),
    .Y(_0751_));
 sky130_fd_sc_hd__o21ai_1 _2102_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[8] ),
    .A2(_0751_),
    .B1(net253),
    .Y(_0752_));
 sky130_fd_sc_hd__nand4_1 _2103_ (.A(_0729_),
    .B(_1044_),
    .C(net37),
    .D(net38),
    .Y(_0753_));
 sky130_fd_sc_hd__a21oi_1 _2104_ (.A1(_0752_),
    .A2(_0753_),
    .B1(_0678_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand4b_4 _2105_ (.A_N(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[10] ),
    .B(net38),
    .C(net37),
    .D(_1044_),
    .Y(_0754_));
 sky130_fd_sc_hd__o31ai_1 _2106_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[9] ),
    .A2(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[8] ),
    .A3(_0746_),
    .B1(net355),
    .Y(_0755_));
 sky130_fd_sc_hd__a21oi_1 _2107_ (.A1(_0754_),
    .A2(_0755_),
    .B1(_0748_),
    .Y(_0251_));
 sky130_fd_sc_hd__o41a_1 _2108_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[10] ),
    .A2(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[9] ),
    .A3(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[8] ),
    .A4(_0746_),
    .B1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .X(_0756_));
 sky130_fd_sc_hd__nor2_1 _2109_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .B(_0754_),
    .Y(_0757_));
 sky130_fd_sc_hd__clkbuf_4 _2110_ (.A(_0684_),
    .X(_0758_));
 sky130_fd_sc_hd__o221a_1 _2111_ (.A1(_1041_),
    .A2(_1046_),
    .B1(_0756_),
    .B2(_0757_),
    .C1(_0758_),
    .X(_0252_));
 sky130_fd_sc_hd__or3_1 _2112_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .C(_0754_),
    .X(_0759_));
 sky130_fd_sc_hd__o21ai_1 _2113_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .A2(_0754_),
    .B1(net373),
    .Y(_0760_));
 sky130_fd_sc_hd__a21oi_1 _2114_ (.A1(_0759_),
    .A2(_0760_),
    .B1(_0748_),
    .Y(_0253_));
 sky130_fd_sc_hd__or4_1 _2115_ (.A(net215),
    .B(_1094_),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[16] ),
    .D(_0746_),
    .X(_0761_));
 sky130_fd_sc_hd__o31a_1 _2116_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ),
    .A2(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .A3(_0754_),
    .B1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[13] ),
    .X(_0762_));
 sky130_fd_sc_hd__nor2_1 _2117_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[13] ),
    .B(_0759_),
    .Y(_0763_));
 sky130_fd_sc_hd__o221a_1 _2118_ (.A1(net219),
    .A2(_0761_),
    .B1(_0762_),
    .B2(_0763_),
    .C1(_0758_),
    .X(_0254_));
 sky130_fd_sc_hd__o41a_1 _2119_ (.A1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[13] ),
    .A2(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ),
    .A3(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .A4(_0754_),
    .B1(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[14] ),
    .X(_0764_));
 sky130_fd_sc_hd__nor4b_1 _2120_ (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ),
    .B(_0754_),
    .C(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ),
    .D_N(_1045_),
    .Y(_0765_));
 sky130_fd_sc_hd__o221a_1 _2121_ (.A1(_1041_),
    .A2(_1046_),
    .B1(_0764_),
    .B2(net33),
    .C1(_0758_),
    .X(_0255_));
 sky130_fd_sc_hd__a21oi_1 _2122_ (.A1(net232),
    .A2(net32),
    .B1(_0748_),
    .Y(_0766_));
 sky130_fd_sc_hd__o21a_1 _2123_ (.A1(net232),
    .A2(net32),
    .B1(_0766_),
    .X(_0256_));
 sky130_fd_sc_hd__or3_1 _2124_ (.A(_1094_),
    .B(net222),
    .C(_0746_),
    .X(_0767_));
 sky130_fd_sc_hd__o21ai_1 _2125_ (.A1(_0746_),
    .A2(_1094_),
    .B1(net222),
    .Y(_0768_));
 sky130_fd_sc_hd__a21oi_1 _2126_ (.A1(_0767_),
    .A2(_0768_),
    .B1(_0748_),
    .Y(_0257_));
 sky130_fd_sc_hd__nand2_1 _2127_ (.A(_0767_),
    .B(net215),
    .Y(_0769_));
 sky130_fd_sc_hd__a21oi_1 _2128_ (.A1(_0761_),
    .A2(_0769_),
    .B1(_0748_),
    .Y(_0258_));
 sky130_fd_sc_hd__o311a_1 _2129_ (.A1(_1042_),
    .A2(_0746_),
    .A3(_1094_),
    .B1(_0721_),
    .C1(net219),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _2130_ (.A(net17),
    .B(_0689_),
    .X(_0770_));
 sky130_fd_sc_hd__clkbuf_1 _2131_ (.A(_0770_),
    .X(_0260_));
 sky130_fd_sc_hd__nor3_2 _2132_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[11] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[10] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ),
    .Y(_0771_));
 sky130_fd_sc_hd__nor3_2 _2133_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[14] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[13] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[12] ),
    .Y(_0772_));
 sky130_fd_sc_hd__inv_2 _2134_ (.A(net372),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_2 _2135_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ),
    .Y(_0774_));
 sky130_fd_sc_hd__nand4_4 _2136_ (.A(_0771_),
    .B(_0772_),
    .C(_0773_),
    .D(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__inv_2 _2137_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[18] ),
    .Y(_0776_));
 sky130_fd_sc_hd__nor2_1 _2138_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[7] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[6] ),
    .Y(_0777_));
 sky130_fd_sc_hd__nor2_1 _2139_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[1] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[0] ),
    .Y(_0778_));
 sky130_fd_sc_hd__nor2_1 _2140_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[3] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[2] ),
    .Y(_0779_));
 sky130_fd_sc_hd__nor2_1 _2141_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[5] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[4] ),
    .Y(_0780_));
 sky130_fd_sc_hd__and4_1 _2142_ (.A(_0777_),
    .B(_0778_),
    .C(_0779_),
    .D(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__buf_2 _2143_ (.A(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__nor2_1 _2144_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[17] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[16] ),
    .Y(_0783_));
 sky130_fd_sc_hd__and4b_1 _2145_ (.A_N(_0775_),
    .B(_0776_),
    .C(_0782_),
    .D(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__clkbuf_4 _2146_ (.A(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__nor3_1 _2147_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[3] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .Y(_0786_));
 sky130_fd_sc_hd__and3_1 _2148_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.rxd_reg ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ),
    .C(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__clkbuf_4 _2149_ (.A(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_4 _2150_ (.A(_0785_),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__nand4_2 _2151_ (.A(_0777_),
    .B(_0778_),
    .C(_0779_),
    .D(_0780_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor4_1 _2152_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[17] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[16] ),
    .C(_0790_),
    .D(_0775_),
    .Y(_0791_));
 sky130_fd_sc_hd__clkbuf_4 _2153_ (.A(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__clkbuf_4 _2154_ (.A(_0776_),
    .X(_0793_));
 sky130_fd_sc_hd__a31o_1 _2155_ (.A1(_0792_),
    .A2(_0788_),
    .A3(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[0] ),
    .X(_0794_));
 sky130_fd_sc_hd__o211a_1 _2156_ (.A1(net208),
    .A2(_0789_),
    .B1(_0794_),
    .C1(_0693_),
    .X(_0261_));
 sky130_fd_sc_hd__a31o_1 _2157_ (.A1(_0792_),
    .A2(_0788_),
    .A3(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[1] ),
    .X(_0795_));
 sky130_fd_sc_hd__o211a_1 _2158_ (.A1(net226),
    .A2(_0789_),
    .B1(_0795_),
    .C1(_0693_),
    .X(_0262_));
 sky130_fd_sc_hd__a31o_1 _2159_ (.A1(_0792_),
    .A2(_0788_),
    .A3(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ),
    .X(_0796_));
 sky130_fd_sc_hd__o211a_1 _2160_ (.A1(net160),
    .A2(_0789_),
    .B1(_0796_),
    .C1(_0693_),
    .X(_0263_));
 sky130_fd_sc_hd__a31o_1 _2161_ (.A1(_0792_),
    .A2(_0788_),
    .A3(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ),
    .X(_0797_));
 sky130_fd_sc_hd__o211a_1 _2162_ (.A1(net221),
    .A2(_0789_),
    .B1(_0797_),
    .C1(_0693_),
    .X(_0264_));
 sky130_fd_sc_hd__a31o_1 _2163_ (.A1(_0792_),
    .A2(_0788_),
    .A3(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[4] ),
    .X(_0798_));
 sky130_fd_sc_hd__o211a_1 _2164_ (.A1(net209),
    .A2(_0789_),
    .B1(_0798_),
    .C1(_0693_),
    .X(_0265_));
 sky130_fd_sc_hd__a31o_1 _2165_ (.A1(_0792_),
    .A2(_0788_),
    .A3(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ),
    .X(_0799_));
 sky130_fd_sc_hd__o211a_1 _2166_ (.A1(net227),
    .A2(_0789_),
    .B1(_0799_),
    .C1(_0693_),
    .X(_0266_));
 sky130_fd_sc_hd__a31o_1 _2167_ (.A1(_0792_),
    .A2(_0788_),
    .A3(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ),
    .X(_0800_));
 sky130_fd_sc_hd__o211a_1 _2168_ (.A1(net234),
    .A2(_0789_),
    .B1(_0800_),
    .C1(_0693_),
    .X(_0267_));
 sky130_fd_sc_hd__a31o_1 _2169_ (.A1(_0792_),
    .A2(_0788_),
    .A3(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[7] ),
    .X(_0801_));
 sky130_fd_sc_hd__o211a_1 _2170_ (.A1(net228),
    .A2(_0789_),
    .B1(_0801_),
    .C1(_0758_),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_4 _2171_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[3] ),
    .X(_0802_));
 sky130_fd_sc_hd__clkbuf_4 _2172_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ),
    .X(_0803_));
 sky130_fd_sc_hd__or2_1 _2173_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ),
    .X(_0804_));
 sky130_fd_sc_hd__clkbuf_4 _2174_ (.A(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__o211ai_2 _2175_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.rxd_reg ),
    .C1(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[3] ),
    .Y(_0806_));
 sky130_fd_sc_hd__o311a_2 _2176_ (.A1(_0802_),
    .A2(_0803_),
    .A3(_0805_),
    .B1(_0806_),
    .C1(_0785_),
    .X(_0807_));
 sky130_fd_sc_hd__nor4_2 _2177_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[3] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .D(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ),
    .Y(_0808_));
 sky130_fd_sc_hd__nand4b_4 _2178_ (.A_N(_0775_),
    .B(_0776_),
    .C(_0782_),
    .D(_0783_),
    .Y(_0809_));
 sky130_fd_sc_hd__a21oi_1 _2179_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.rxd_reg ),
    .A2(_0808_),
    .B1(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _2180_ (.A(net369),
    .B(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__o211a_1 _2181_ (.A1(net369),
    .A2(_0807_),
    .B1(_0811_),
    .C1(_0758_),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_1 _2182_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ),
    .Y(_0812_));
 sky130_fd_sc_hd__nand2_1 _2183_ (.A(_0805_),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__a221o_1 _2184_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.rxd_reg ),
    .A2(_0808_),
    .B1(_0806_),
    .B2(_0813_),
    .C1(_0809_),
    .X(_0814_));
 sky130_fd_sc_hd__o211a_1 _2185_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .A2(_0810_),
    .B1(_0721_),
    .C1(_0814_),
    .X(_0270_));
 sky130_fd_sc_hd__and3_2 _2186_ (.A(net31),
    .B(_0806_),
    .C(_0776_),
    .X(_0815_));
 sky130_fd_sc_hd__nor4b_1 _2187_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ),
    .D_N(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[3] ),
    .Y(_0816_));
 sky130_fd_sc_hd__a21o_1 _2188_ (.A1(_0805_),
    .A2(_0803_),
    .B1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__a22oi_1 _2189_ (.A1(_0803_),
    .A2(_0809_),
    .B1(_0815_),
    .B2(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_1 _2190_ (.A(_0678_),
    .B(_0818_),
    .Y(_0271_));
 sky130_fd_sc_hd__o31a_1 _2191_ (.A1(_0803_),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .A3(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ),
    .B1(_0802_),
    .X(_0819_));
 sky130_fd_sc_hd__o211ai_1 _2192_ (.A1(_0808_),
    .A2(_0819_),
    .B1(_0806_),
    .C1(_0810_),
    .Y(_0820_));
 sky130_fd_sc_hd__nand2_1 _2193_ (.A(_0809_),
    .B(_0802_),
    .Y(_0821_));
 sky130_fd_sc_hd__a21oi_1 _2194_ (.A1(_0820_),
    .A2(_0821_),
    .B1(_0678_),
    .Y(_0272_));
 sky130_fd_sc_hd__clkbuf_4 _2195_ (.A(_0809_),
    .X(_0822_));
 sky130_fd_sc_hd__o21ai_1 _2196_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.rxd_reg ),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ),
    .B1(_0786_),
    .Y(_0823_));
 sky130_fd_sc_hd__clkbuf_4 _2197_ (.A(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__a21oi_1 _2198_ (.A1(_0792_),
    .A2(_0793_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[0] ),
    .Y(_0825_));
 sky130_fd_sc_hd__o221a_1 _2199_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0825_),
    .B2(_0807_),
    .C1(_0758_),
    .X(_0273_));
 sky130_fd_sc_hd__and2_1 _2200_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[1] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[0] ),
    .X(_0826_));
 sky130_fd_sc_hd__o2bb2a_1 _2201_ (.A1_N(_0776_),
    .A2_N(net31),
    .B1(_0826_),
    .B2(_0778_),
    .X(_0827_));
 sky130_fd_sc_hd__o221a_1 _2202_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0827_),
    .B2(_0815_),
    .C1(_0758_),
    .X(_0274_));
 sky130_fd_sc_hd__o21a_1 _2203_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[1] ),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[0] ),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[2] ),
    .X(_0828_));
 sky130_fd_sc_hd__nor3_1 _2204_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[2] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[1] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[0] ),
    .Y(_0829_));
 sky130_fd_sc_hd__o2bb2a_1 _2205_ (.A1_N(_0776_),
    .A2_N(net31),
    .B1(_0828_),
    .B2(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__o221a_1 _2206_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0830_),
    .B2(_0815_),
    .C1(_0758_),
    .X(_0275_));
 sky130_fd_sc_hd__nand2_1 _2207_ (.A(_0778_),
    .B(_0779_),
    .Y(_0831_));
 sky130_fd_sc_hd__o31ai_1 _2208_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[2] ),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[1] ),
    .A3(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[0] ),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[3] ),
    .Y(_0832_));
 sky130_fd_sc_hd__a21oi_1 _2209_ (.A1(_0831_),
    .A2(_0832_),
    .B1(_0785_),
    .Y(_0833_));
 sky130_fd_sc_hd__o221a_1 _2210_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0833_),
    .B2(_0815_),
    .C1(_0758_),
    .X(_0276_));
 sky130_fd_sc_hd__or4b_1 _2211_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[4] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[3] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[2] ),
    .D_N(_0778_),
    .X(_0834_));
 sky130_fd_sc_hd__nand2_1 _2212_ (.A(_0831_),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[4] ),
    .Y(_0835_));
 sky130_fd_sc_hd__a21oi_1 _2213_ (.A1(_0834_),
    .A2(_0835_),
    .B1(_0785_),
    .Y(_0836_));
 sky130_fd_sc_hd__o221a_1 _2214_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0836_),
    .B2(_0807_),
    .C1(_0721_),
    .X(_0277_));
 sky130_fd_sc_hd__or3_1 _2215_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[5] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[4] ),
    .C(_0831_),
    .X(_0837_));
 sky130_fd_sc_hd__o21ai_1 _2216_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[4] ),
    .A2(_0831_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[5] ),
    .Y(_0838_));
 sky130_fd_sc_hd__a21oi_1 _2217_ (.A1(_0837_),
    .A2(_0838_),
    .B1(_0785_),
    .Y(_0839_));
 sky130_fd_sc_hd__and3_1 _2218_ (.A(net31),
    .B(_0808_),
    .C(_0776_),
    .X(_0840_));
 sky130_fd_sc_hd__o221a_1 _2219_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0839_),
    .B2(_0840_),
    .C1(_0721_),
    .X(_0278_));
 sky130_fd_sc_hd__nand2_1 _2220_ (.A(_0837_),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[6] ),
    .Y(_0841_));
 sky130_fd_sc_hd__or4_1 _2221_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[6] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[5] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[4] ),
    .D(_0831_),
    .X(_0842_));
 sky130_fd_sc_hd__a21oi_1 _2222_ (.A1(_0841_),
    .A2(_0842_),
    .B1(_0785_),
    .Y(_0843_));
 sky130_fd_sc_hd__o221a_1 _2223_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0843_),
    .B2(_0807_),
    .C1(_0721_),
    .X(_0279_));
 sky130_fd_sc_hd__buf_2 _2224_ (.A(_0790_),
    .X(_0844_));
 sky130_fd_sc_hd__nand2_1 _2225_ (.A(_0842_),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[7] ),
    .Y(_0845_));
 sky130_fd_sc_hd__a21oi_1 _2226_ (.A1(_0844_),
    .A2(_0845_),
    .B1(_0785_),
    .Y(_0846_));
 sky130_fd_sc_hd__o21a_1 _2227_ (.A1(_0809_),
    .A2(_0824_),
    .B1(_0684_),
    .X(_0847_));
 sky130_fd_sc_hd__o21a_1 _2228_ (.A1(_0840_),
    .A2(_0846_),
    .B1(_0847_),
    .X(_0280_));
 sky130_fd_sc_hd__nand2_1 _2229_ (.A(_0844_),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ),
    .Y(_0848_));
 sky130_fd_sc_hd__nand2_1 _2230_ (.A(_0782_),
    .B(_0774_),
    .Y(_0849_));
 sky130_fd_sc_hd__a21oi_1 _2231_ (.A1(_0848_),
    .A2(_0849_),
    .B1(_0785_),
    .Y(_0850_));
 sky130_fd_sc_hd__o221a_1 _2232_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0850_),
    .B2(_0815_),
    .C1(_0721_),
    .X(_0281_));
 sky130_fd_sc_hd__o21ai_1 _2233_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ),
    .A2(_0844_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ),
    .Y(_0851_));
 sky130_fd_sc_hd__or3_1 _2234_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ),
    .C(_0844_),
    .X(_0852_));
 sky130_fd_sc_hd__a21oi_1 _2235_ (.A1(_0851_),
    .A2(_0852_),
    .B1(_0785_),
    .Y(_0853_));
 sky130_fd_sc_hd__o221a_1 _2236_ (.A1(_0809_),
    .A2(_0824_),
    .B1(_0853_),
    .B2(_0807_),
    .C1(_0721_),
    .X(_0282_));
 sky130_fd_sc_hd__or4_1 _2237_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[10] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ),
    .D(_0790_),
    .X(_0854_));
 sky130_fd_sc_hd__o21ai_1 _2238_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ),
    .A2(_0849_),
    .B1(net264),
    .Y(_0855_));
 sky130_fd_sc_hd__a21o_1 _2239_ (.A1(net31),
    .A2(_0793_),
    .B1(_0677_),
    .X(_0856_));
 sky130_fd_sc_hd__a21oi_1 _2240_ (.A1(_0854_),
    .A2(_0855_),
    .B1(_0856_),
    .Y(_0283_));
 sky130_fd_sc_hd__or3_1 _2241_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[16] ),
    .B(_0844_),
    .C(_0775_),
    .X(_0857_));
 sky130_fd_sc_hd__a32o_1 _2242_ (.A1(_0774_),
    .A2(_0782_),
    .A3(_0771_),
    .B1(_0854_),
    .B2(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[11] ),
    .X(_0858_));
 sky130_fd_sc_hd__o311a_1 _2243_ (.A1(net212),
    .A2(net328),
    .A3(_0857_),
    .B1(_0684_),
    .C1(_0858_),
    .X(_0284_));
 sky130_fd_sc_hd__or4_2 _2244_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[11] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[10] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ),
    .D(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ),
    .X(_0859_));
 sky130_fd_sc_hd__o41a_1 _2245_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[7] ),
    .A2(_0859_),
    .A3(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[6] ),
    .A4(_0837_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[12] ),
    .X(_0860_));
 sky130_fd_sc_hd__and4b_1 _2246_ (.A_N(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[12] ),
    .B(_0782_),
    .C(_0771_),
    .D(_0774_),
    .X(_0861_));
 sky130_fd_sc_hd__o211a_1 _2247_ (.A1(_0860_),
    .A2(_0861_),
    .B1(_0721_),
    .C1(_0822_),
    .X(_0285_));
 sky130_fd_sc_hd__or4_1 _2248_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[13] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[12] ),
    .C(_0844_),
    .D(_0859_),
    .X(_0862_));
 sky130_fd_sc_hd__o31ai_1 _2249_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[12] ),
    .A2(_0844_),
    .A3(_0859_),
    .B1(net220),
    .Y(_0863_));
 sky130_fd_sc_hd__a21oi_1 _2250_ (.A1(_0862_),
    .A2(_0863_),
    .B1(_0856_),
    .Y(_0286_));
 sky130_fd_sc_hd__nor4_1 _2251_ (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[11] ),
    .B(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[10] ),
    .C(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ),
    .D(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ),
    .Y(_0864_));
 sky130_fd_sc_hd__a32oi_1 _2252_ (.A1(_0782_),
    .A2(net36),
    .A3(_0772_),
    .B1(_0862_),
    .B2(net211),
    .Y(_0865_));
 sky130_fd_sc_hd__nor2_1 _2253_ (.A(_0856_),
    .B(_0865_),
    .Y(_0287_));
 sky130_fd_sc_hd__or4b_1 _2254_ (.A(net372),
    .B(_0844_),
    .C(_0859_),
    .D_N(_0772_),
    .X(_0866_));
 sky130_fd_sc_hd__a31o_1 _2255_ (.A1(_0782_),
    .A2(_0864_),
    .A3(_0772_),
    .B1(_0773_),
    .X(_0867_));
 sky130_fd_sc_hd__a21oi_1 _2256_ (.A1(_0866_),
    .A2(_0867_),
    .B1(_0856_),
    .Y(_0288_));
 sky130_fd_sc_hd__o21ai_1 _2257_ (.A1(_0844_),
    .A2(_0775_),
    .B1(net367),
    .Y(_0868_));
 sky130_fd_sc_hd__a21oi_1 _2258_ (.A1(_0857_),
    .A2(_0868_),
    .B1(_0856_),
    .Y(_0289_));
 sky130_fd_sc_hd__o31a_1 _2259_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[16] ),
    .A2(_0844_),
    .A3(_0775_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[17] ),
    .X(_0869_));
 sky130_fd_sc_hd__o211a_1 _2260_ (.A1(_0792_),
    .A2(_0869_),
    .B1(_0822_),
    .C1(_0758_),
    .X(_0290_));
 sky130_fd_sc_hd__o311a_1 _2261_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[17] ),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[16] ),
    .A3(_0866_),
    .B1(_0684_),
    .C1(net212),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_4 _2262_ (.A(_0627_),
    .X(_0870_));
 sky130_fd_sc_hd__clkbuf_4 _2263_ (.A(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__nand3_4 _2264_ (.A(_0643_),
    .B(_0660_),
    .C(_0593_),
    .Y(_0872_));
 sky130_fd_sc_hd__a32o_1 _2265_ (.A1(_0587_),
    .A2(_0871_),
    .A3(_0661_),
    .B1(_0872_),
    .B2(net81),
    .X(_0292_));
 sky130_fd_sc_hd__a32o_1 _2266_ (.A1(_0597_),
    .A2(_0871_),
    .A3(_0661_),
    .B1(_0872_),
    .B2(net96),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_4 _2267_ (.A(_0660_),
    .X(_0873_));
 sky130_fd_sc_hd__a32o_1 _2268_ (.A1(_0489_),
    .A2(_0871_),
    .A3(_0873_),
    .B1(_0872_),
    .B2(net80),
    .X(_0294_));
 sky130_fd_sc_hd__a32o_1 _2269_ (.A1(_0491_),
    .A2(_0871_),
    .A3(_0873_),
    .B1(_0872_),
    .B2(net111),
    .X(_0295_));
 sky130_fd_sc_hd__a32o_1 _2270_ (.A1(_0601_),
    .A2(_0871_),
    .A3(_0873_),
    .B1(_0872_),
    .B2(net83),
    .X(_0296_));
 sky130_fd_sc_hd__a32o_1 _2271_ (.A1(_0494_),
    .A2(_0871_),
    .A3(_0873_),
    .B1(_0872_),
    .B2(net101),
    .X(_0297_));
 sky130_fd_sc_hd__a32o_1 _2272_ (.A1(_0496_),
    .A2(_0871_),
    .A3(_0873_),
    .B1(_0872_),
    .B2(net107),
    .X(_0298_));
 sky130_fd_sc_hd__a32o_1 _2273_ (.A1(_0605_),
    .A2(_0870_),
    .A3(_0873_),
    .B1(_0872_),
    .B2(net93),
    .X(_0299_));
 sky130_fd_sc_hd__nand3_4 _2274_ (.A(_0643_),
    .B(_0479_),
    .C(_0660_),
    .Y(_0874_));
 sky130_fd_sc_hd__a32o_1 _2275_ (.A1(_0587_),
    .A2(_0710_),
    .A3(_0873_),
    .B1(_0874_),
    .B2(net128),
    .X(_0300_));
 sky130_fd_sc_hd__a32o_1 _2276_ (.A1(_0597_),
    .A2(_0710_),
    .A3(_0873_),
    .B1(_0874_),
    .B2(net122),
    .X(_0301_));
 sky130_fd_sc_hd__a32o_1 _2277_ (.A1(_0489_),
    .A2(_0710_),
    .A3(_0873_),
    .B1(_0874_),
    .B2(net138),
    .X(_0302_));
 sky130_fd_sc_hd__a32o_1 _2278_ (.A1(_0491_),
    .A2(_0710_),
    .A3(_0873_),
    .B1(_0874_),
    .B2(net114),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_4 _2279_ (.A(_0660_),
    .X(_0875_));
 sky130_fd_sc_hd__a32o_1 _2280_ (.A1(_0601_),
    .A2(_0710_),
    .A3(_0875_),
    .B1(_0874_),
    .B2(net157),
    .X(_0304_));
 sky130_fd_sc_hd__a32o_1 _2281_ (.A1(_0494_),
    .A2(_0710_),
    .A3(_0875_),
    .B1(_0874_),
    .B2(net94),
    .X(_0305_));
 sky130_fd_sc_hd__a32o_1 _2282_ (.A1(_0496_),
    .A2(_0486_),
    .A3(_0875_),
    .B1(_0874_),
    .B2(net146),
    .X(_0306_));
 sky130_fd_sc_hd__a32o_1 _2283_ (.A1(_0605_),
    .A2(_0486_),
    .A3(_0875_),
    .B1(_0874_),
    .B2(net102),
    .X(_0307_));
 sky130_fd_sc_hd__o2111ai_4 _2284_ (.A1(_0589_),
    .A2(_0590_),
    .B1(_0592_),
    .C1(_0627_),
    .D1(_0972_),
    .Y(_0876_));
 sky130_fd_sc_hd__a22o_1 _2285_ (.A1(_0876_),
    .A2(net193),
    .B1(_0484_),
    .B2(_0871_),
    .X(_0308_));
 sky130_fd_sc_hd__a22o_1 _2286_ (.A1(_0876_),
    .A2(net188),
    .B1(_0488_),
    .B2(_0871_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2287_ (.A0(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ),
    .A1(net269),
    .S(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__clkbuf_1 _2288_ (.A(_0877_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2289_ (.A0(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ),
    .A1(net271),
    .S(_0876_),
    .X(_0878_));
 sky130_fd_sc_hd__clkbuf_1 _2290_ (.A(_0878_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2291_ (.A0(_0601_),
    .A1(net306),
    .S(_0876_),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_1 _2292_ (.A(_0879_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2293_ (.A0(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ),
    .A1(net267),
    .S(_0876_),
    .X(_0880_));
 sky130_fd_sc_hd__clkbuf_1 _2294_ (.A(_0880_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2295_ (.A0(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ),
    .A1(net284),
    .S(_0876_),
    .X(_0881_));
 sky130_fd_sc_hd__clkbuf_1 _2296_ (.A(_0881_),
    .X(_0314_));
 sky130_fd_sc_hd__a22o_1 _2297_ (.A1(_0876_),
    .A2(net158),
    .B1(_0498_),
    .B2(_0871_),
    .X(_0315_));
 sky130_fd_sc_hd__nand3_4 _2298_ (.A(_0643_),
    .B(_0641_),
    .C(_0593_),
    .Y(_0882_));
 sky130_fd_sc_hd__a32o_1 _2299_ (.A1(_0587_),
    .A2(_0870_),
    .A3(_0709_),
    .B1(_0882_),
    .B2(net109),
    .X(_0316_));
 sky130_fd_sc_hd__a32o_1 _2300_ (.A1(_0597_),
    .A2(_0870_),
    .A3(_0709_),
    .B1(_0882_),
    .B2(net95),
    .X(_0317_));
 sky130_fd_sc_hd__a32o_1 _2301_ (.A1(_0489_),
    .A2(_0870_),
    .A3(_0709_),
    .B1(_0882_),
    .B2(net92),
    .X(_0318_));
 sky130_fd_sc_hd__a32o_1 _2302_ (.A1(_0491_),
    .A2(_0870_),
    .A3(_0709_),
    .B1(_0882_),
    .B2(net91),
    .X(_0319_));
 sky130_fd_sc_hd__a32o_1 _2303_ (.A1(_0601_),
    .A2(_0870_),
    .A3(_0673_),
    .B1(_0882_),
    .B2(net112),
    .X(_0320_));
 sky130_fd_sc_hd__a32o_1 _2304_ (.A1(_0494_),
    .A2(_0870_),
    .A3(_0673_),
    .B1(_0882_),
    .B2(net124),
    .X(_0321_));
 sky130_fd_sc_hd__a32o_1 _2305_ (.A1(_0496_),
    .A2(_0870_),
    .A3(_0673_),
    .B1(_0882_),
    .B2(net90),
    .X(_0322_));
 sky130_fd_sc_hd__a32o_1 _2306_ (.A1(_0605_),
    .A2(_0870_),
    .A3(_0673_),
    .B1(_0882_),
    .B2(net108),
    .X(_0323_));
 sky130_fd_sc_hd__nand4_1 _2307_ (.A(net370),
    .B(_0476_),
    .C(_0975_),
    .D(_0980_),
    .Y(_0883_));
 sky130_fd_sc_hd__a21oi_1 _2308_ (.A1(_0789_),
    .A2(_0883_),
    .B1(_0678_),
    .Y(_0324_));
 sky130_fd_sc_hd__nand3b_4 _2309_ (.A_N(_0643_),
    .B(_0660_),
    .C(_0593_),
    .Y(_0884_));
 sky130_fd_sc_hd__a32o_1 _2310_ (.A1(_0587_),
    .A2(_0875_),
    .A3(_0666_),
    .B1(_0884_),
    .B2(net99),
    .X(_0325_));
 sky130_fd_sc_hd__a32o_1 _2311_ (.A1(_0597_),
    .A2(_0875_),
    .A3(_0666_),
    .B1(_0884_),
    .B2(net127),
    .X(_0326_));
 sky130_fd_sc_hd__a32o_1 _2312_ (.A1(_0489_),
    .A2(_0875_),
    .A3(_0666_),
    .B1(_0884_),
    .B2(net97),
    .X(_0327_));
 sky130_fd_sc_hd__a32o_1 _2313_ (.A1(_0491_),
    .A2(_0875_),
    .A3(_0666_),
    .B1(_0884_),
    .B2(net72),
    .X(_0328_));
 sky130_fd_sc_hd__a32o_1 _2314_ (.A1(_0601_),
    .A2(_0875_),
    .A3(_0666_),
    .B1(_0884_),
    .B2(net79),
    .X(_0329_));
 sky130_fd_sc_hd__a32o_1 _2315_ (.A1(_0494_),
    .A2(_0875_),
    .A3(_0666_),
    .B1(_0884_),
    .B2(net104),
    .X(_0330_));
 sky130_fd_sc_hd__a32o_1 _2316_ (.A1(_0496_),
    .A2(_0660_),
    .A3(_0666_),
    .B1(_0884_),
    .B2(net106),
    .X(_0331_));
 sky130_fd_sc_hd__a32o_1 _2317_ (.A1(_0605_),
    .A2(_0660_),
    .A3(_0666_),
    .B1(_0884_),
    .B2(net85),
    .X(_0332_));
 sky130_fd_sc_hd__o31a_1 _2318_ (.A1(_0802_),
    .A2(_0803_),
    .A3(_0805_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[1] ),
    .X(_0885_));
 sky130_fd_sc_hd__o21ai_1 _2319_ (.A1(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[3] ),
    .Y(_0886_));
 sky130_fd_sc_hd__nand3_1 _2320_ (.A(_0823_),
    .B(net6),
    .C(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__nor2_4 _2321_ (.A(_0809_),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(net208),
    .A1(_0885_),
    .S(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_1 _2323_ (.A(_0889_),
    .X(_0333_));
 sky130_fd_sc_hd__o31a_1 _2324_ (.A1(_0802_),
    .A2(_0803_),
    .A3(_0805_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[2] ),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _2325_ (.A0(net226),
    .A1(_0890_),
    .S(_0888_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_1 _2326_ (.A(_0891_),
    .X(_0334_));
 sky130_fd_sc_hd__o31a_1 _2327_ (.A1(_0802_),
    .A2(_0803_),
    .A3(_0805_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[3] ),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _2328_ (.A0(net160),
    .A1(_0892_),
    .S(_0888_),
    .X(_0893_));
 sky130_fd_sc_hd__clkbuf_1 _2329_ (.A(_0893_),
    .X(_0335_));
 sky130_fd_sc_hd__o31a_1 _2330_ (.A1(_0802_),
    .A2(_0803_),
    .A3(_0805_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[4] ),
    .X(_0894_));
 sky130_fd_sc_hd__mux2_1 _2331_ (.A0(net221),
    .A1(_0894_),
    .S(_0888_),
    .X(_0895_));
 sky130_fd_sc_hd__clkbuf_1 _2332_ (.A(_0895_),
    .X(_0336_));
 sky130_fd_sc_hd__o31a_1 _2333_ (.A1(_0802_),
    .A2(_0803_),
    .A3(_0805_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[5] ),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(net209),
    .A1(_0896_),
    .S(_0888_),
    .X(_0897_));
 sky130_fd_sc_hd__clkbuf_1 _2335_ (.A(_0897_),
    .X(_0337_));
 sky130_fd_sc_hd__o31a_1 _2336_ (.A1(_0802_),
    .A2(_0803_),
    .A3(_0805_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[6] ),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _2337_ (.A0(net227),
    .A1(_0898_),
    .S(_0888_),
    .X(_0899_));
 sky130_fd_sc_hd__clkbuf_1 _2338_ (.A(_0899_),
    .X(_0338_));
 sky130_fd_sc_hd__o31a_1 _2339_ (.A1(_0802_),
    .A2(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ),
    .A3(_0805_),
    .B1(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[7] ),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _2340_ (.A0(net234),
    .A1(_0900_),
    .S(_0888_),
    .X(_0901_));
 sky130_fd_sc_hd__clkbuf_1 _2341_ (.A(_0901_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(net228),
    .A1(\uart_inst.uart_core_inst.uart_rx_inst.rxd_reg ),
    .S(_0888_),
    .X(_0902_));
 sky130_fd_sc_hd__clkbuf_1 _2343_ (.A(_0902_),
    .X(_0340_));
 sky130_fd_sc_hd__o311a_2 _2344_ (.A1(_0934_),
    .A2(_0401_),
    .A3(_0465_),
    .B1(\uart_inst.uart_core_inst.uart_tx_inst.s_axis_tready_reg ),
    .C1(_1052_),
    .X(_0903_));
 sky130_fd_sc_hd__a21oi_1 _2345_ (.A1(_1090_),
    .A2(net310),
    .B1(_1052_),
    .Y(_0904_));
 sky130_fd_sc_hd__nor3_1 _2346_ (.A(_0903_),
    .B(_0678_),
    .C(_0904_),
    .Y(_0341_));
 sky130_fd_sc_hd__o21ai_1 _2347_ (.A1(_1080_),
    .A2(_0903_),
    .B1(_0684_),
    .Y(_0905_));
 sky130_fd_sc_hd__a21oi_1 _2348_ (.A1(_1080_),
    .A2(_0903_),
    .B1(_0905_),
    .Y(_0342_));
 sky130_fd_sc_hd__and2_1 _2349_ (.A(_1077_),
    .B(\uart_inst.uart_core_inst.uart_tx_inst.s_axis_tready_reg ),
    .X(_0906_));
 sky130_fd_sc_hd__a31o_1 _2350_ (.A1(_1090_),
    .A2(_0906_),
    .A3(_1080_),
    .B1(_1064_),
    .X(_0907_));
 sky130_fd_sc_hd__o2111ai_2 _2351_ (.A1(_0403_),
    .A2(_0719_),
    .B1(_0906_),
    .C1(_1080_),
    .D1(_1064_),
    .Y(_0908_));
 sky130_fd_sc_hd__and3_1 _2352_ (.A(_0907_),
    .B(_0908_),
    .C(_1037_),
    .X(_0909_));
 sky130_fd_sc_hd__clkbuf_1 _2353_ (.A(_0909_),
    .X(_0343_));
 sky130_fd_sc_hd__nor2_1 _2354_ (.A(_1087_),
    .B(_0925_),
    .Y(_0910_));
 sky130_fd_sc_hd__a31o_1 _2355_ (.A1(_1080_),
    .A2(_0903_),
    .A3(_0910_),
    .B1(_0677_),
    .X(_0911_));
 sky130_fd_sc_hd__a21oi_1 _2356_ (.A1(_1087_),
    .A2(_0908_),
    .B1(_0911_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand4_1 _2357_ (.A(\uart_inst.fifo_tx_inst.read_ptr_reg[4] ),
    .B(_1080_),
    .C(_0903_),
    .D(_0910_),
    .Y(_0912_));
 sky130_fd_sc_hd__a41o_1 _2358_ (.A1(_1090_),
    .A2(_0906_),
    .A3(_0910_),
    .A4(_1080_),
    .B1(\uart_inst.fifo_tx_inst.read_ptr_reg[4] ),
    .X(_0913_));
 sky130_fd_sc_hd__and3_1 _2359_ (.A(_0912_),
    .B(_0913_),
    .C(_1037_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_1 _2360_ (.A(_0914_),
    .X(_0345_));
 sky130_fd_sc_hd__a21oi_1 _2361_ (.A1(_0544_),
    .A2(_0473_),
    .B1(_0689_),
    .Y(_0915_));
 sky130_fd_sc_hd__o21a_1 _2362_ (.A1(_0544_),
    .A2(_0473_),
    .B1(_0915_),
    .X(_0346_));
 sky130_fd_sc_hd__a21o_1 _2363_ (.A1(_0416_),
    .A2(_0444_),
    .B1(_0440_),
    .X(_0916_));
 sky130_fd_sc_hd__and3_1 _2364_ (.A(_0916_),
    .B(_1037_),
    .C(_0504_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_1 _2365_ (.A(_0917_),
    .X(_0347_));
 sky130_fd_sc_hd__a21oi_1 _2366_ (.A1(_0558_),
    .A2(_0502_),
    .B1(_0689_),
    .Y(_0918_));
 sky130_fd_sc_hd__o21a_1 _2367_ (.A1(_0558_),
    .A2(_0502_),
    .B1(_0918_),
    .X(_0348_));
 sky130_fd_sc_hd__and4_1 _2368_ (.A(_0506_),
    .B(_0443_),
    .C(_0439_),
    .D(_0545_),
    .X(_0919_));
 sky130_fd_sc_hd__a21boi_1 _2369_ (.A1(_0558_),
    .A2(_0502_),
    .B1_N(_0451_),
    .Y(_0920_));
 sky130_fd_sc_hd__o21a_1 _2370_ (.A1(_0919_),
    .A2(_0920_),
    .B1(_0693_),
    .X(_0349_));
 sky130_fd_sc_hd__nand4_1 _2371_ (.A(\uart_inst.fifo_tx_inst.write_ptr_reg[4] ),
    .B(_0451_),
    .C(_0412_),
    .D(_0501_),
    .Y(_0921_));
 sky130_fd_sc_hd__and3_1 _2372_ (.A(_0413_),
    .B(_0412_),
    .C(_0928_),
    .X(_0922_));
 sky130_fd_sc_hd__a31o_1 _2373_ (.A1(_0440_),
    .A2(_0438_),
    .A3(_0922_),
    .B1(\uart_inst.fifo_tx_inst.write_ptr_reg[4] ),
    .X(_0923_));
 sky130_fd_sc_hd__and3_1 _2374_ (.A(_0921_),
    .B(_1037_),
    .C(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__clkbuf_1 _2375_ (.A(_0924_),
    .X(_0350_));
 sky130_fd_sc_hd__dfxtp_1 _2376_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0000_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2377_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0001_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2378_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0002_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2379_ (.CLK(clknet_leaf_22_PCLK),
    .D(net176),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2380_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0004_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2381_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0005_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2382_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0006_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2383_ (.CLK(clknet_leaf_13_PCLK),
    .D(net150),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2384_ (.CLK(clknet_leaf_11_PCLK),
    .D(_0008_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2385_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0009_),
    .Q(\uart_inst.fifo_tx_inst.mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2386_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0010_),
    .Q(\uart_inst.fifo_tx_inst.mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2387_ (.CLK(clknet_leaf_25_PCLK),
    .D(_0011_),
    .Q(\uart_inst.fifo_tx_inst.mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2388_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0012_),
    .Q(\uart_inst.fifo_tx_inst.mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2389_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0013_),
    .Q(\uart_inst.fifo_tx_inst.mem[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2390_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0014_),
    .Q(\uart_inst.fifo_tx_inst.mem[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2391_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0015_),
    .Q(\uart_inst.fifo_tx_inst.mem[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2392_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0016_),
    .Q(\uart_inst.fifo_tx_inst.mem[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2393_ (.CLK(clknet_leaf_25_PCLK),
    .D(_0017_),
    .Q(\uart_inst.fifo_tx_inst.mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2394_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0018_),
    .Q(\uart_inst.fifo_tx_inst.mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2395_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0019_),
    .Q(\uart_inst.fifo_tx_inst.mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2396_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0020_),
    .Q(\uart_inst.fifo_tx_inst.mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2397_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0021_),
    .Q(\uart_inst.fifo_tx_inst.mem[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2398_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0022_),
    .Q(\uart_inst.fifo_tx_inst.mem[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2399_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0023_),
    .Q(\uart_inst.fifo_tx_inst.mem[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2400_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0024_),
    .Q(\uart_inst.fifo_tx_inst.mem[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2401_ (.CLK(clknet_leaf_25_PCLK),
    .D(_0025_),
    .Q(\uart_inst.fifo_tx_inst.mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2402_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0026_),
    .Q(\uart_inst.fifo_tx_inst.mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2403_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0027_),
    .Q(\uart_inst.fifo_tx_inst.mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2404_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0028_),
    .Q(\uart_inst.fifo_tx_inst.mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2405_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0029_),
    .Q(\uart_inst.fifo_tx_inst.mem[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2406_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0030_),
    .Q(\uart_inst.fifo_tx_inst.mem[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2407_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0031_),
    .Q(\uart_inst.fifo_tx_inst.mem[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2408_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0032_),
    .Q(\uart_inst.fifo_tx_inst.mem[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2409_ (.CLK(clknet_leaf_25_PCLK),
    .D(_0033_),
    .Q(\uart_inst.fifo_tx_inst.mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2410_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0034_),
    .Q(\uart_inst.fifo_tx_inst.mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2411_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0035_),
    .Q(\uart_inst.fifo_tx_inst.mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2412_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0036_),
    .Q(\uart_inst.fifo_tx_inst.mem[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2413_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0037_),
    .Q(\uart_inst.fifo_tx_inst.mem[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2414_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0038_),
    .Q(\uart_inst.fifo_tx_inst.mem[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2415_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0039_),
    .Q(\uart_inst.fifo_tx_inst.mem[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2416_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0040_),
    .Q(\uart_inst.fifo_tx_inst.mem[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2417_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0041_),
    .Q(\uart_inst.fifo_rx_inst.mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2418_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0042_),
    .Q(\uart_inst.fifo_rx_inst.mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2419_ (.CLK(clknet_leaf_1_PCLK),
    .D(_0043_),
    .Q(\uart_inst.fifo_rx_inst.mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2420_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0044_),
    .Q(\uart_inst.fifo_rx_inst.mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2421_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0045_),
    .Q(\uart_inst.fifo_rx_inst.mem[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2422_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0046_),
    .Q(\uart_inst.fifo_rx_inst.mem[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2423_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0047_),
    .Q(\uart_inst.fifo_rx_inst.mem[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2424_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0048_),
    .Q(\uart_inst.fifo_rx_inst.mem[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2425_ (.CLK(clknet_leaf_20_PCLK),
    .D(_0049_),
    .Q(\uart_inst.fifo_tx_inst.mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2426_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0050_),
    .Q(\uart_inst.fifo_tx_inst.mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2427_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0051_),
    .Q(\uart_inst.fifo_tx_inst.mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2428_ (.CLK(clknet_leaf_20_PCLK),
    .D(_0052_),
    .Q(\uart_inst.fifo_tx_inst.mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2429_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0053_),
    .Q(\uart_inst.fifo_tx_inst.mem[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2430_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0054_),
    .Q(\uart_inst.fifo_tx_inst.mem[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2431_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0055_),
    .Q(\uart_inst.fifo_tx_inst.mem[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2432_ (.CLK(clknet_leaf_20_PCLK),
    .D(_0056_),
    .Q(\uart_inst.fifo_tx_inst.mem[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2433_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0057_),
    .Q(\uart_inst.fifo_tx_inst.mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2434_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0058_),
    .Q(\uart_inst.fifo_tx_inst.mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2435_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0059_),
    .Q(\uart_inst.fifo_tx_inst.mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2436_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0060_),
    .Q(\uart_inst.fifo_tx_inst.mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2437_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0061_),
    .Q(\uart_inst.fifo_tx_inst.mem[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2438_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0062_),
    .Q(\uart_inst.fifo_tx_inst.mem[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2439_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0063_),
    .Q(\uart_inst.fifo_tx_inst.mem[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2440_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0064_),
    .Q(\uart_inst.fifo_tx_inst.mem[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2441_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0065_),
    .Q(\uart_inst.fifo_tx_inst.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2442_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0066_),
    .Q(\uart_inst.fifo_tx_inst.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2443_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0067_),
    .Q(\uart_inst.fifo_tx_inst.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2444_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0068_),
    .Q(\uart_inst.fifo_tx_inst.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2445_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0069_),
    .Q(\uart_inst.fifo_tx_inst.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2446_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0070_),
    .Q(\uart_inst.fifo_tx_inst.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2447_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0071_),
    .Q(\uart_inst.fifo_tx_inst.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2448_ (.CLK(clknet_leaf_14_PCLK),
    .D(_0072_),
    .Q(\uart_inst.fifo_tx_inst.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2449_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0073_),
    .Q(\uart_inst.fifo_tx_inst.mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2450_ (.CLK(clknet_leaf_25_PCLK),
    .D(_0074_),
    .Q(\uart_inst.fifo_tx_inst.mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2451_ (.CLK(clknet_leaf_25_PCLK),
    .D(_0075_),
    .Q(\uart_inst.fifo_tx_inst.mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2452_ (.CLK(clknet_leaf_25_PCLK),
    .D(_0076_),
    .Q(\uart_inst.fifo_tx_inst.mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2453_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0077_),
    .Q(\uart_inst.fifo_tx_inst.mem[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2454_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0078_),
    .Q(\uart_inst.fifo_tx_inst.mem[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2455_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0079_),
    .Q(\uart_inst.fifo_tx_inst.mem[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2456_ (.CLK(clknet_leaf_17_PCLK),
    .D(_0080_),
    .Q(\uart_inst.fifo_tx_inst.mem[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2457_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0081_),
    .Q(\uart_inst.fifo_tx_inst.mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2458_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0082_),
    .Q(\uart_inst.fifo_tx_inst.mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2459_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0083_),
    .Q(\uart_inst.fifo_tx_inst.mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2460_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0084_),
    .Q(\uart_inst.fifo_tx_inst.mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2461_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0085_),
    .Q(\uart_inst.fifo_tx_inst.mem[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2462_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0086_),
    .Q(\uart_inst.fifo_tx_inst.mem[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2463_ (.CLK(clknet_leaf_21_PCLK),
    .D(_0087_),
    .Q(\uart_inst.fifo_tx_inst.mem[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2464_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0088_),
    .Q(\uart_inst.fifo_tx_inst.mem[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2465_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0089_),
    .Q(\uart_inst.fifo_tx_inst.mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2466_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0090_),
    .Q(\uart_inst.fifo_tx_inst.mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2467_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0091_),
    .Q(\uart_inst.fifo_tx_inst.mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2468_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0092_),
    .Q(\uart_inst.fifo_tx_inst.mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2469_ (.CLK(clknet_leaf_21_PCLK),
    .D(_0093_),
    .Q(\uart_inst.fifo_tx_inst.mem[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2470_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0094_),
    .Q(\uart_inst.fifo_tx_inst.mem[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2471_ (.CLK(clknet_leaf_20_PCLK),
    .D(_0095_),
    .Q(\uart_inst.fifo_tx_inst.mem[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2472_ (.CLK(clknet_leaf_21_PCLK),
    .D(_0096_),
    .Q(\uart_inst.fifo_tx_inst.mem[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2473_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0097_),
    .Q(\uart_inst.fifo_tx_inst.mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2474_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0098_),
    .Q(\uart_inst.fifo_tx_inst.mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2475_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0099_),
    .Q(\uart_inst.fifo_tx_inst.mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2476_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0100_),
    .Q(\uart_inst.fifo_tx_inst.mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2477_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0101_),
    .Q(\uart_inst.fifo_tx_inst.mem[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2478_ (.CLK(clknet_leaf_14_PCLK),
    .D(_0102_),
    .Q(\uart_inst.fifo_tx_inst.mem[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2479_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0103_),
    .Q(\uart_inst.fifo_tx_inst.mem[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2480_ (.CLK(clknet_leaf_14_PCLK),
    .D(_0104_),
    .Q(\uart_inst.fifo_tx_inst.mem[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2481_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0105_),
    .Q(\uart_inst.fifo_tx_inst.mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2482_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0106_),
    .Q(\uart_inst.fifo_tx_inst.mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2483_ (.CLK(clknet_leaf_21_PCLK),
    .D(_0107_),
    .Q(\uart_inst.fifo_tx_inst.mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2484_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0108_),
    .Q(\uart_inst.fifo_tx_inst.mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2485_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0109_),
    .Q(\uart_inst.fifo_tx_inst.mem[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2486_ (.CLK(clknet_leaf_14_PCLK),
    .D(_0110_),
    .Q(\uart_inst.fifo_tx_inst.mem[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2487_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0111_),
    .Q(\uart_inst.fifo_tx_inst.mem[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2488_ (.CLK(clknet_leaf_14_PCLK),
    .D(_0112_),
    .Q(\uart_inst.fifo_tx_inst.mem[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2489_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0113_),
    .Q(\uart_inst.fifo_tx_inst.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2490_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0114_),
    .Q(\uart_inst.fifo_tx_inst.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2491_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0115_),
    .Q(\uart_inst.fifo_tx_inst.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2492_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0116_),
    .Q(\uart_inst.fifo_tx_inst.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2493_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0117_),
    .Q(\uart_inst.fifo_tx_inst.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2494_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0118_),
    .Q(\uart_inst.fifo_tx_inst.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2495_ (.CLK(clknet_leaf_20_PCLK),
    .D(_0119_),
    .Q(\uart_inst.fifo_tx_inst.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2496_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0120_),
    .Q(\uart_inst.fifo_tx_inst.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2497_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0121_),
    .Q(\uart_inst.fifo_rx_inst.mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2498_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0122_),
    .Q(\uart_inst.fifo_rx_inst.mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2499_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0123_),
    .Q(\uart_inst.fifo_rx_inst.mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2500_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0124_),
    .Q(\uart_inst.fifo_rx_inst.mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2501_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0125_),
    .Q(\uart_inst.fifo_rx_inst.mem[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2502_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0126_),
    .Q(\uart_inst.fifo_rx_inst.mem[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2503_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0127_),
    .Q(\uart_inst.fifo_rx_inst.mem[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2504_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0128_),
    .Q(\uart_inst.fifo_rx_inst.mem[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2505_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0129_),
    .Q(\uart_inst.fifo_tx_inst.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2506_ (.CLK(clknet_leaf_23_PCLK),
    .D(_0130_),
    .Q(\uart_inst.fifo_tx_inst.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2507_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0131_),
    .Q(\uart_inst.fifo_tx_inst.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2508_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0132_),
    .Q(\uart_inst.fifo_tx_inst.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2509_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0133_),
    .Q(\uart_inst.fifo_tx_inst.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2510_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0134_),
    .Q(\uart_inst.fifo_tx_inst.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2511_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0135_),
    .Q(\uart_inst.fifo_tx_inst.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2512_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0136_),
    .Q(\uart_inst.fifo_tx_inst.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2513_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0137_),
    .Q(\uart_inst.fifo_tx_inst.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2514_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0138_),
    .Q(\uart_inst.fifo_tx_inst.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2515_ (.CLK(clknet_leaf_27_PCLK),
    .D(_0139_),
    .Q(\uart_inst.fifo_tx_inst.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2516_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0140_),
    .Q(\uart_inst.fifo_tx_inst.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2517_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0141_),
    .Q(\uart_inst.fifo_tx_inst.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2518_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0142_),
    .Q(\uart_inst.fifo_tx_inst.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2519_ (.CLK(clknet_leaf_16_PCLK),
    .D(_0143_),
    .Q(\uart_inst.fifo_tx_inst.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2520_ (.CLK(clknet_leaf_15_PCLK),
    .D(_0144_),
    .Q(\uart_inst.fifo_tx_inst.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2521_ (.CLK(clknet_leaf_25_PCLK),
    .D(_0145_),
    .Q(\uart_inst.fifo_tx_inst.mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2522_ (.CLK(clknet_leaf_24_PCLK),
    .D(_0146_),
    .Q(\uart_inst.fifo_tx_inst.mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2523_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0147_),
    .Q(\uart_inst.fifo_tx_inst.mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2524_ (.CLK(clknet_leaf_26_PCLK),
    .D(_0148_),
    .Q(\uart_inst.fifo_tx_inst.mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2525_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0149_),
    .Q(\uart_inst.fifo_tx_inst.mem[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2526_ (.CLK(clknet_leaf_18_PCLK),
    .D(_0150_),
    .Q(\uart_inst.fifo_tx_inst.mem[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2527_ (.CLK(clknet_leaf_19_PCLK),
    .D(_0151_),
    .Q(\uart_inst.fifo_tx_inst.mem[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2528_ (.CLK(clknet_leaf_20_PCLK),
    .D(_0152_),
    .Q(\uart_inst.fifo_tx_inst.mem[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2529_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0153_),
    .Q(\uart_inst.fifo_rx_inst.mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2530_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0154_),
    .Q(\uart_inst.fifo_rx_inst.mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2531_ (.CLK(clknet_leaf_1_PCLK),
    .D(_0155_),
    .Q(\uart_inst.fifo_rx_inst.mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2532_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0156_),
    .Q(\uart_inst.fifo_rx_inst.mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2533_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0157_),
    .Q(\uart_inst.fifo_rx_inst.mem[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2534_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0158_),
    .Q(\uart_inst.fifo_rx_inst.mem[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2535_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0159_),
    .Q(\uart_inst.fifo_rx_inst.mem[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2536_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0160_),
    .Q(\uart_inst.fifo_rx_inst.mem[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2537_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0161_),
    .Q(\uart_inst.fifo_rx_inst.mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2538_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0162_),
    .Q(\uart_inst.fifo_rx_inst.mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2539_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0163_),
    .Q(\uart_inst.fifo_rx_inst.mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2540_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0164_),
    .Q(\uart_inst.fifo_rx_inst.mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2541_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0165_),
    .Q(\uart_inst.fifo_rx_inst.mem[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2542_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0166_),
    .Q(\uart_inst.fifo_rx_inst.mem[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2543_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0167_),
    .Q(\uart_inst.fifo_rx_inst.mem[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2544_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0168_),
    .Q(\uart_inst.fifo_rx_inst.mem[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2545_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0169_),
    .Q(\uart_inst.fifo_rx_inst.mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2546_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0170_),
    .Q(\uart_inst.fifo_rx_inst.mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2547_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0171_),
    .Q(\uart_inst.fifo_rx_inst.mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2548_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0172_),
    .Q(\uart_inst.fifo_rx_inst.mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2549_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0173_),
    .Q(\uart_inst.fifo_rx_inst.mem[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2550_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0174_),
    .Q(\uart_inst.fifo_rx_inst.mem[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2551_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0175_),
    .Q(\uart_inst.fifo_rx_inst.mem[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2552_ (.CLK(clknet_leaf_27_PCLK),
    .D(_0176_),
    .Q(\uart_inst.fifo_rx_inst.mem[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2553_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0177_),
    .Q(\uart_inst.fifo_rx_inst.mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2554_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0178_),
    .Q(\uart_inst.fifo_rx_inst.mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2555_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0179_),
    .Q(\uart_inst.fifo_rx_inst.mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2556_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0180_),
    .Q(\uart_inst.fifo_rx_inst.mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2557_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0181_),
    .Q(\uart_inst.fifo_rx_inst.mem[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2558_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0182_),
    .Q(\uart_inst.fifo_rx_inst.mem[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2559_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0183_),
    .Q(\uart_inst.fifo_rx_inst.mem[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2560_ (.CLK(clknet_leaf_27_PCLK),
    .D(_0184_),
    .Q(\uart_inst.fifo_rx_inst.mem[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2561_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0185_),
    .Q(\uart_inst.fifo_rx_inst.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2562_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0186_),
    .Q(\uart_inst.fifo_rx_inst.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2563_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0187_),
    .Q(\uart_inst.fifo_rx_inst.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2564_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0188_),
    .Q(\uart_inst.fifo_rx_inst.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2565_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0189_),
    .Q(\uart_inst.fifo_rx_inst.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2566_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0190_),
    .Q(\uart_inst.fifo_rx_inst.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2567_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0191_),
    .Q(\uart_inst.fifo_rx_inst.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2568_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0192_),
    .Q(\uart_inst.fifo_rx_inst.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2569_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0193_),
    .Q(\uart_inst.fifo_rx_inst.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2570_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0194_),
    .Q(\uart_inst.fifo_rx_inst.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2571_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0195_),
    .Q(\uart_inst.fifo_rx_inst.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2572_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0196_),
    .Q(\uart_inst.fifo_rx_inst.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2573_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0197_),
    .Q(\uart_inst.fifo_rx_inst.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2574_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0198_),
    .Q(\uart_inst.fifo_rx_inst.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2575_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0199_),
    .Q(\uart_inst.fifo_rx_inst.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2576_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0200_),
    .Q(\uart_inst.fifo_rx_inst.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2577_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0201_),
    .Q(\uart_inst.fifo_rx_inst.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2578_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0202_),
    .Q(\uart_inst.fifo_rx_inst.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2579_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0203_),
    .Q(\uart_inst.fifo_rx_inst.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2580_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0204_),
    .Q(\uart_inst.fifo_rx_inst.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2581_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0205_),
    .Q(\uart_inst.fifo_rx_inst.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2582_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0206_),
    .Q(\uart_inst.fifo_rx_inst.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2583_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0207_),
    .Q(\uart_inst.fifo_rx_inst.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2584_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0208_),
    .Q(\uart_inst.fifo_rx_inst.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2585_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0209_),
    .Q(\uart_inst.fifo_rx_inst.read_ptr_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2586_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0210_),
    .Q(\uart_inst.fifo_rx_inst.read_ptr_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2587_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0211_),
    .Q(\uart_inst.fifo_rx_inst.read_ptr_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2588_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0212_),
    .Q(\uart_inst.fifo_rx_inst.read_ptr_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2589_ (.CLK(clknet_leaf_12_PCLK),
    .D(_0213_),
    .Q(\uart_inst.fifo_rx_inst.read_ptr_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2590_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0214_),
    .Q(\uart_inst.fifo_rx_inst.write_ptr_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2591_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0215_),
    .Q(\uart_inst.fifo_rx_inst.write_ptr_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2592_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0216_),
    .Q(\uart_inst.fifo_rx_inst.write_ptr_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2593_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0217_),
    .Q(\uart_inst.fifo_rx_inst.write_ptr_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2594_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0218_),
    .Q(\uart_inst.fifo_rx_inst.write_ptr_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2595_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0219_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _2596_ (.CLK(clknet_leaf_11_PCLK),
    .D(_0220_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.s_axis_tready_reg ));
 sky130_fd_sc_hd__dfxtp_1 _2597_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0221_),
    .Q(\uart_inst.fifo_rx_inst.mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2598_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0222_),
    .Q(\uart_inst.fifo_rx_inst.mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2599_ (.CLK(clknet_leaf_1_PCLK),
    .D(_0223_),
    .Q(\uart_inst.fifo_rx_inst.mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2600_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0224_),
    .Q(\uart_inst.fifo_rx_inst.mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2601_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0225_),
    .Q(\uart_inst.fifo_rx_inst.mem[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2602_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0226_),
    .Q(\uart_inst.fifo_rx_inst.mem[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2603_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0227_),
    .Q(\uart_inst.fifo_rx_inst.mem[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2604_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0228_),
    .Q(\uart_inst.fifo_rx_inst.mem[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2605_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0229_),
    .Q(\uart_inst.fifo_rx_inst.mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2606_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0230_),
    .Q(\uart_inst.fifo_rx_inst.mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2607_ (.CLK(clknet_leaf_1_PCLK),
    .D(_0231_),
    .Q(\uart_inst.fifo_rx_inst.mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2608_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0232_),
    .Q(\uart_inst.fifo_rx_inst.mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2609_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0233_),
    .Q(\uart_inst.fifo_rx_inst.mem[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2610_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0234_),
    .Q(\uart_inst.fifo_rx_inst.mem[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2611_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0235_),
    .Q(\uart_inst.fifo_rx_inst.mem[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2612_ (.CLK(clknet_leaf_31_PCLK),
    .D(_0236_),
    .Q(\uart_inst.fifo_rx_inst.mem[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2613_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0237_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2614_ (.CLK(clknet_leaf_11_PCLK),
    .D(net334),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2615_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0239_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2616_ (.CLK(clknet_leaf_3_PCLK),
    .D(_0240_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2617_ (.CLK(clknet_leaf_10_PCLK),
    .D(_0241_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2618_ (.CLK(clknet_leaf_14_PCLK),
    .D(_0242_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2619_ (.CLK(clknet_leaf_14_PCLK),
    .D(_0243_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2620_ (.CLK(clknet_leaf_10_PCLK),
    .D(_0244_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2621_ (.CLK(clknet_leaf_10_PCLK),
    .D(_0245_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2622_ (.CLK(clknet_leaf_10_PCLK),
    .D(_0246_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2623_ (.CLK(clknet_leaf_14_PCLK),
    .D(net218),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2624_ (.CLK(clknet_leaf_10_PCLK),
    .D(_0248_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2625_ (.CLK(clknet_leaf_11_PCLK),
    .D(_0249_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2626_ (.CLK(clknet_leaf_11_PCLK),
    .D(_0250_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2627_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0251_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _2628_ (.CLK(clknet_leaf_11_PCLK),
    .D(_0252_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2629_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0253_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2630_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0254_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2631_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0255_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2632_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0256_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2633_ (.CLK(clknet_leaf_10_PCLK),
    .D(_0257_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2634_ (.CLK(clknet_leaf_9_PCLK),
    .D(net216),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2635_ (.CLK(clknet_leaf_11_PCLK),
    .D(_0259_),
    .Q(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _2636_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0260_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.rxd_reg ));
 sky130_fd_sc_hd__dfxtp_1 _2637_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0261_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2638_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0262_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2639_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0263_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[2] ));
 sky130_fd_sc_hd__dfxtp_4 _2640_ (.CLK(clknet_leaf_5_PCLK),
    .D(_0264_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2641_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0265_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2642_ (.CLK(clknet_leaf_5_PCLK),
    .D(_0266_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2643_ (.CLK(clknet_leaf_5_PCLK),
    .D(_0267_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2644_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0268_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tdata_reg[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2645_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0269_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2646_ (.CLK(clknet_leaf_11_PCLK),
    .D(_0270_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2647_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0271_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2648_ (.CLK(clknet_leaf_11_PCLK),
    .D(_0272_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2649_ (.CLK(clknet_leaf_6_PCLK),
    .D(_0273_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2650_ (.CLK(clknet_leaf_7_PCLK),
    .D(_0274_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2651_ (.CLK(clknet_leaf_7_PCLK),
    .D(_0275_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2652_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0276_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2653_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0277_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2654_ (.CLK(clknet_leaf_9_PCLK),
    .D(_0278_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2655_ (.CLK(clknet_leaf_8_PCLK),
    .D(_0279_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2656_ (.CLK(clknet_leaf_7_PCLK),
    .D(_0280_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2657_ (.CLK(clknet_leaf_7_PCLK),
    .D(_0281_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2658_ (.CLK(clknet_leaf_7_PCLK),
    .D(_0282_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2659_ (.CLK(clknet_leaf_7_PCLK),
    .D(_0283_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2660_ (.CLK(clknet_leaf_6_PCLK),
    .D(_0284_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2661_ (.CLK(clknet_leaf_8_PCLK),
    .D(_0285_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2662_ (.CLK(clknet_leaf_8_PCLK),
    .D(_0286_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2663_ (.CLK(clknet_leaf_8_PCLK),
    .D(_0287_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2664_ (.CLK(clknet_leaf_6_PCLK),
    .D(_0288_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2665_ (.CLK(clknet_leaf_6_PCLK),
    .D(_0289_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2666_ (.CLK(clknet_leaf_6_PCLK),
    .D(_0290_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2667_ (.CLK(clknet_leaf_6_PCLK),
    .D(net213),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2668_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0292_),
    .Q(\uart_inst.fifo_rx_inst.mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2669_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0293_),
    .Q(\uart_inst.fifo_rx_inst.mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2670_ (.CLK(clknet_leaf_1_PCLK),
    .D(_0294_),
    .Q(\uart_inst.fifo_rx_inst.mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2671_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0295_),
    .Q(\uart_inst.fifo_rx_inst.mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2672_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0296_),
    .Q(\uart_inst.fifo_rx_inst.mem[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2673_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0297_),
    .Q(\uart_inst.fifo_rx_inst.mem[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2674_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0298_),
    .Q(\uart_inst.fifo_rx_inst.mem[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2675_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0299_),
    .Q(\uart_inst.fifo_rx_inst.mem[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2676_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0300_),
    .Q(\uart_inst.fifo_rx_inst.mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2677_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0301_),
    .Q(\uart_inst.fifo_rx_inst.mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2678_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0302_),
    .Q(\uart_inst.fifo_rx_inst.mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2679_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0303_),
    .Q(\uart_inst.fifo_rx_inst.mem[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2680_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0304_),
    .Q(\uart_inst.fifo_rx_inst.mem[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2681_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0305_),
    .Q(\uart_inst.fifo_rx_inst.mem[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2682_ (.CLK(clknet_leaf_0_PCLK),
    .D(_0306_),
    .Q(\uart_inst.fifo_rx_inst.mem[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2683_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0307_),
    .Q(\uart_inst.fifo_rx_inst.mem[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2684_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0308_),
    .Q(\uart_inst.fifo_rx_inst.mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2685_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0309_),
    .Q(\uart_inst.fifo_rx_inst.mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2686_ (.CLK(clknet_leaf_1_PCLK),
    .D(_0310_),
    .Q(\uart_inst.fifo_rx_inst.mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2687_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0311_),
    .Q(\uart_inst.fifo_rx_inst.mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2688_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0312_),
    .Q(\uart_inst.fifo_rx_inst.mem[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2689_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0313_),
    .Q(\uart_inst.fifo_rx_inst.mem[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2690_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0314_),
    .Q(\uart_inst.fifo_rx_inst.mem[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2691_ (.CLK(clknet_leaf_33_PCLK),
    .D(_0315_),
    .Q(\uart_inst.fifo_rx_inst.mem[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2692_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0316_),
    .Q(\uart_inst.fifo_rx_inst.mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2693_ (.CLK(clknet_leaf_2_PCLK),
    .D(_0317_),
    .Q(\uart_inst.fifo_rx_inst.mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2694_ (.CLK(clknet_leaf_1_PCLK),
    .D(_0318_),
    .Q(\uart_inst.fifo_rx_inst.mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2695_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0319_),
    .Q(\uart_inst.fifo_rx_inst.mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2696_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0320_),
    .Q(\uart_inst.fifo_rx_inst.mem[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2697_ (.CLK(clknet_leaf_36_PCLK),
    .D(_0321_),
    .Q(\uart_inst.fifo_rx_inst.mem[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2698_ (.CLK(clknet_leaf_35_PCLK),
    .D(_0322_),
    .Q(\uart_inst.fifo_rx_inst.mem[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2699_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0323_),
    .Q(\uart_inst.fifo_rx_inst.mem[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2700_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0324_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tvalid_reg ));
 sky130_fd_sc_hd__dfxtp_1 _2701_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0325_),
    .Q(\uart_inst.fifo_rx_inst.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2702_ (.CLK(clknet_leaf_30_PCLK),
    .D(_0326_),
    .Q(\uart_inst.fifo_rx_inst.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2703_ (.CLK(clknet_leaf_29_PCLK),
    .D(_0327_),
    .Q(\uart_inst.fifo_rx_inst.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2704_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0328_),
    .Q(\uart_inst.fifo_rx_inst.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2705_ (.CLK(clknet_leaf_28_PCLK),
    .D(_0329_),
    .Q(\uart_inst.fifo_rx_inst.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2706_ (.CLK(clknet_leaf_34_PCLK),
    .D(_0330_),
    .Q(\uart_inst.fifo_rx_inst.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2707_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0331_),
    .Q(\uart_inst.fifo_rx_inst.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2708_ (.CLK(clknet_leaf_32_PCLK),
    .D(_0332_),
    .Q(\uart_inst.fifo_rx_inst.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2709_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0333_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2710_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0334_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2711_ (.CLK(clknet_leaf_5_PCLK),
    .D(_0335_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2712_ (.CLK(clknet_leaf_5_PCLK),
    .D(_0336_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2713_ (.CLK(clknet_leaf_5_PCLK),
    .D(_0337_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2714_ (.CLK(clknet_leaf_5_PCLK),
    .D(_0338_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2715_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0339_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2716_ (.CLK(clknet_leaf_4_PCLK),
    .D(_0340_),
    .Q(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2717_ (.CLK(clknet_leaf_12_PCLK),
    .D(_0341_),
    .Q(\uart_inst.fifo_tx_inst.read_ptr_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2718_ (.CLK(clknet_leaf_12_PCLK),
    .D(_0342_),
    .Q(\uart_inst.fifo_tx_inst.read_ptr_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2719_ (.CLK(clknet_leaf_12_PCLK),
    .D(_0343_),
    .Q(\uart_inst.fifo_tx_inst.read_ptr_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2720_ (.CLK(clknet_leaf_12_PCLK),
    .D(_0344_),
    .Q(\uart_inst.fifo_tx_inst.read_ptr_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2721_ (.CLK(clknet_leaf_12_PCLK),
    .D(_0345_),
    .Q(\uart_inst.fifo_tx_inst.read_ptr_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2722_ (.CLK(clknet_leaf_12_PCLK),
    .D(_0346_),
    .Q(\uart_inst.fifo_tx_inst.write_ptr_reg[0] ));
 sky130_fd_sc_hd__dfxtp_4 _2723_ (.CLK(clknet_leaf_12_PCLK),
    .D(_0347_),
    .Q(\uart_inst.fifo_tx_inst.write_ptr_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2724_ (.CLK(clknet_leaf_13_PCLK),
    .D(_0348_),
    .Q(\uart_inst.fifo_tx_inst.write_ptr_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2725_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0349_),
    .Q(\uart_inst.fifo_tx_inst.write_ptr_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2726_ (.CLK(clknet_leaf_22_PCLK),
    .D(_0350_),
    .Q(\uart_inst.fifo_tx_inst.write_ptr_reg[4] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_PCLK (.A(PCLK),
    .X(clknet_0_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_PCLK (.A(clknet_0_PCLK),
    .X(clknet_2_0__leaf_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_PCLK (.A(clknet_0_PCLK),
    .X(clknet_2_1__leaf_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_PCLK (.A(clknet_0_PCLK),
    .X(clknet_2_2__leaf_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_PCLK (.A(clknet_0_PCLK),
    .X(clknet_2_3__leaf_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_0_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_10_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_11_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_12_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_13_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_14_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_15_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_16_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_17_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_18_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_19_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_1_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_20_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_PCLK (.A(clknet_2_3__leaf_PCLK),
    .X(clknet_leaf_21_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_22_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_23_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_24_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_25_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_26_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_27_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_28_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_29_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_2_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_PCLK (.A(clknet_2_2__leaf_PCLK),
    .X(clknet_leaf_30_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_31_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_32_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_33_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_34_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_35_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_PCLK (.A(clknet_2_0__leaf_PCLK),
    .X(clknet_leaf_36_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_3_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_4_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_5_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_6_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_7_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_8_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_PCLK (.A(clknet_2_1__leaf_PCLK),
    .X(clknet_leaf_9_PCLK));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\uart_inst.fifo_rx_inst.mem[4][7] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\uart_inst.fifo_rx_inst.mem[4][1] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\uart_inst.fifo_rx_inst.mem[6][0] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\uart_inst.fifo_rx_inst.mem[6][1] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\uart_inst.fifo_tx_inst.mem[11][1] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\uart_inst.fifo_tx_inst.mem[14][1] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\uart_inst.fifo_tx_inst.mem[11][2] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\uart_inst.fifo_tx_inst.mem[15][2] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\uart_inst.fifo_tx_inst.mem[10][7] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\uart_inst.fifo_tx_inst.mem[3][3] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[3] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0003_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\uart_inst.fifo_rx_inst.mem[14][3] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\uart_inst.fifo_rx_inst.mem[3][0] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\uart_inst.fifo_rx_inst.mem[3][2] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\uart_inst.fifo_rx_inst.mem[3][4] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[2] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\uart_inst.fifo_rx_inst.mem[3][7] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\uart_inst.fifo_tx_inst.mem[6][1] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\uart_inst.fifo_rx_inst.mem[1][1] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\uart_inst.fifo_rx_inst.mem[5][2] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\uart_inst.fifo_rx_inst.mem[1][0] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[1] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\uart_inst.fifo_rx_inst.mem[0][4] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\uart_inst.fifo_rx_inst.mem[13][4] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\uart_inst.fifo_rx_inst.mem[11][1] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\uart_inst.fifo_tx_inst.mem[10][3] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\uart_inst.fifo_rx_inst.mem[1][7] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\uart_inst.fifo_rx_inst.mem[1][4] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[8] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\uart_inst.fifo_rx_inst.mem[11][0] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\uart_inst.fifo_tx_inst.mem[15][0] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\uart_inst.fifo_tx_inst.mem[3][2] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\uart_inst.fifo_tx_inst.mem[11][5] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\uart_inst.fifo_rx_inst.mem[8][2] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\uart_inst.fifo_tx_inst.mem[11][6] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\uart_inst.fifo_tx_inst.mem[3][0] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\uart_inst.fifo_tx_inst.mem[2][1] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\uart_inst.fifo_tx_inst.mem[6][3] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\uart_inst.fifo_rx_inst.mem[3][1] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\uart_inst.fifo_tx_inst.mem[6][6] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\uart_inst.fifo_tx_inst.mem[6][7] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[7] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0747_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\uart_inst.fifo_tx_inst.mem[11][4] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\uart_inst.fifo_rx_inst.mem[8][0] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[0] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[0] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[4] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\uart_inst.fifo_tx_inst.mem[15][4] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[14] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[18] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0291_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[4] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[17] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0258_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\uart_inst.fifo_rx_inst.mem[2][3] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[6] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0247_),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[18] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[13] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[3] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[16] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\uart_inst.fifo_tx_inst.mem[7][1] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\uart_inst.fifo_tx_inst.mem[7][2] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\uart_inst.fifo_tx_inst.mem[3][5] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[1] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\uart_inst.fifo_rx_inst.mem[8][4] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[5] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[7] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\uart_inst.fifo_tx_inst.mem[11][0] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\uart_inst.fifo_tx_inst.mem[3][6] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\uart_inst.fifo_tx_inst.mem[3][4] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[15] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\uart_inst.fifo_tx_inst.mem[7][4] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[6] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\uart_inst.fifo_tx_inst.mem[11][7] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\uart_inst.fifo_tx_inst.mem[3][7] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\uart_inst.fifo_rx_inst.mem[6][3] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\uart_inst.fifo_tx_inst.mem[7][6] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\uart_inst.fifo_tx_inst.mem[7][3] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\uart_inst.fifo_tx_inst.mem[7][0] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\uart_inst.fifo_tx_inst.mem[15][7] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\uart_inst.fifo_tx_inst.mem[11][3] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\uart_inst.fifo_rx_inst.mem[13][2] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\uart_inst.fifo_tx_inst.mem[7][7] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\uart_inst.fifo_rx_inst.mem[9][2] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\uart_inst.fifo_rx_inst.mem[7][7] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\uart_inst.fifo_rx_inst.mem[9][0] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\uart_inst.fifo_rx_inst.mem[0][7] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\uart_inst.fifo_tx_inst.mem[10][4] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\uart_inst.fifo_tx_inst.mem[7][5] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\uart_inst.fifo_rx_inst.mem[9][6] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\uart_inst.fifo_rx_inst.mem[7][1] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\uart_inst.fifo_rx_inst.mem[9][1] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\uart_inst.fifo_rx_inst.mem[7][5] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[9] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\uart_inst.fifo_tx_inst.mem[10][6] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\uart_inst.fifo_rx_inst.mem[7][3] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\uart_inst.fifo_rx_inst.mem[9][5] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\uart_inst.fifo_rx_inst.mem[4][3] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\uart_inst.fifo_tx_inst.mem[12][6] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\uart_inst.fifo_tx_inst.mem[12][7] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\uart_inst.fifo_rx_inst.mem[9][4] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\uart_inst.fifo_rx_inst.mem[13][1] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\uart_inst.fifo_rx_inst.mem[7][0] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\uart_inst.fifo_rx_inst.mem[9][7] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\uart_inst.fifo_tx_inst.mem[10][1] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[10] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\uart_inst.fifo_tx_inst.mem[10][2] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\uart_inst.fifo_rx_inst.mem[7][6] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\uart_inst.fifo_rx_inst.mem[6][7] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\uart_inst.fifo_rx_inst.mem[4][4] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\uart_inst.fifo_rx_inst.mem[11][5] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\uart_inst.fifo_rx_inst.mem[13][6] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\uart_inst.fifo_rx_inst.mem[11][2] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\uart_inst.fifo_tx_inst.mem[5][1] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\uart_inst.fifo_rx_inst.mem[11][3] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\uart_inst.fifo_tx_inst.mem[8][4] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\uart_inst.fifo_rx_inst.mem[7][2] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\uart_inst.fifo_rx_inst.mem[15][2] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\uart_inst.fifo_tx_inst.mem[13][6] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\uart_inst.fifo_tx_inst.mem[2][3] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\uart_inst.fifo_rx_inst.mem[4][6] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\uart_inst.fifo_tx_inst.mem[0][3] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\uart_inst.fifo_rx_inst.mem[7][4] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\uart_inst.fifo_tx_inst.mem[13][2] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\uart_inst.fifo_rx_inst.mem[13][3] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\uart_inst.fifo_tx_inst.mem[12][2] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\uart_inst.fifo_tx_inst.mem[2][0] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\uart_inst.fifo_rx_inst.mem[15][6] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\uart_inst.fifo_rx_inst.mem[11][6] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\uart_inst.fifo_rx_inst.mem[13][0] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\uart_inst.fifo_tx_inst.mem[2][6] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\uart_inst.fifo_rx_inst.mem[6][6] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\uart_inst.fifo_tx_inst.mem[13][1] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\uart_inst.fifo_rx_inst.mem[9][3] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\uart_inst.fifo_tx_inst.mem[13][7] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\uart_inst.fifo_tx_inst.mem[13][0] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\uart_inst.fifo_tx_inst.mem[12][3] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\uart_inst.fifo_tx_inst.mem[5][2] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\uart_inst.fifo_tx_inst.mem[4][6] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\uart_inst.fifo_tx_inst.mem[9][5] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\uart_inst.fifo_tx_inst.mem[13][4] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\uart_inst.fifo_tx_inst.mem[5][7] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\uart_inst.fifo_rx_inst.mem[10][6] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\uart_inst.fifo_tx_inst.mem[14][4] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\uart_inst.fifo_tx_inst.mem[4][5] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\uart_inst.fifo_rx_inst.mem[15][3] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\uart_inst.fifo_tx_inst.mem[13][3] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\uart_inst.fifo_tx_inst.mem[8][7] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\uart_inst.fifo_tx_inst.mem[9][7] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\uart_inst.fifo_tx_inst.mem[1][3] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\uart_inst.fifo_tx_inst.mem[4][0] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\uart_inst.fifo_tx_inst.mem[5][4] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\uart_inst.fifo_rx_inst.mem[11][4] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\uart_inst.fifo_rx_inst.mem[10][3] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\uart_inst.fifo_tx_inst.mem[0][7] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\uart_inst.fifo_tx_inst.mem[4][1] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\uart_inst.fifo_tx_inst.mem[8][1] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\uart_inst.uart_core_inst.uart_tx_inst.s_axis_tready_reg ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\uart_inst.fifo_tx_inst.mem[5][3] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\uart_inst.fifo_tx_inst.mem[12][0] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\uart_inst.fifo_tx_inst.mem[14][0] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\uart_inst.fifo_rx_inst.mem[15][5] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\uart_inst.fifo_tx_inst.mem[14][2] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\uart_inst.fifo_tx_inst.mem[9][0] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\uart_inst.fifo_rx_inst.mem[10][2] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\uart_inst.fifo_tx_inst.mem[8][5] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\uart_inst.fifo_tx_inst.mem[12][1] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\uart_inst.fifo_tx_inst.mem[9][4] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\uart_inst.fifo_tx_inst.mem[0][0] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\uart_inst.fifo_tx_inst.mem[3][1] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\uart_inst.fifo_tx_inst.mem[5][6] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\uart_inst.fifo_tx_inst.mem[9][1] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\uart_inst.fifo_tx_inst.mem[0][5] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\uart_inst.fifo_tx_inst.mem[13][5] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\uart_inst.fifo_tx_inst.mem[8][2] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\uart_inst.fifo_rx_inst.mem[8][7] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\uart_inst.fifo_rx_inst.mem[13][5] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[17] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\uart_inst.fifo_tx_inst.mem[8][0] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\uart_inst.fifo_tx_inst.mem[1][0] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\uart_inst.fifo_tx_inst.mem[4][7] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[5] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[1] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0238_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\uart_inst.fifo_tx_inst.mem[14][3] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\uart_inst.fifo_tx_inst.mem[9][2] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\uart_inst.fifo_rx_inst.mem[12][5] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[1] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\uart_inst.fifo_tx_inst.mem[6][0] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\uart_inst.fifo_tx_inst.mem[6][5] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\uart_inst.fifo_tx_inst.mem[12][4] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\uart_inst.fifo_tx_inst.mem[9][3] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\uart_inst.fifo_tx_inst.mem[8][3] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\uart_inst.fifo_tx_inst.mem[5][5] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\uart_inst.fifo_tx_inst.mem[2][2] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\uart_inst.fifo_tx_inst.mem[4][3] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\uart_inst.fifo_tx_inst.mem[8][6] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\uart_inst.fifo_rx_inst.mem[10][1] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\uart_inst.fifo_tx_inst.mem[1][1] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\uart_inst.fifo_tx_inst.mem[9][6] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\uart_inst.fifo_tx_inst.mem[0][4] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\uart_inst.fifo_tx_inst.mem[0][1] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\uart_inst.uart_core_inst.uart_tx_inst.bit_cnt[3] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\uart_inst.fifo_tx_inst.mem[0][6] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\uart_inst.fifo_tx_inst.mem[10][5] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\uart_inst.fifo_tx_inst.mem[2][5] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[10] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net26),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\uart_inst.fifo_rx_inst.mem[8][1] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\uart_inst.fifo_rx_inst.read_ptr_reg[4] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\uart_inst.fifo_tx_inst.mem[1][2] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\uart_inst.fifo_tx_inst.mem[1][6] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\uart_inst.fifo_tx_inst.mem[10][0] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\uart_inst.fifo_tx_inst.mem[2][7] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\uart_inst.fifo_tx_inst.mem[2][4] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\uart_inst.fifo_tx_inst.mem[0][2] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\uart_inst.fifo_tx_inst.mem[1][5] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\uart_inst.fifo_tx_inst.mem[1][4] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\uart_inst.fifo_tx_inst.mem[5][0] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\uart_inst.fifo_rx_inst.mem[14][2] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\uart_inst.fifo_rx_inst.mem[0][2] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[16] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\uart_inst.fifo_tx_inst.mem[1][7] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\uart_inst.uart_core_inst.uart_rx_inst.bit_cnt[0] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\uart_inst.uart_core_inst.uart_rx_inst.m_axis_tvalid_reg ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[8] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\uart_inst.uart_core_inst.uart_rx_inst.prescale_reg[15] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\uart_inst.uart_core_inst.uart_tx_inst.prescale_reg[12] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\uart_inst.fifo_rx_inst.write_ptr_reg[0] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\uart_inst.fifo_rx_inst.mem[2][2] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\uart_inst.fifo_rx_inst.mem[0][0] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\uart_inst.fifo_rx_inst.mem[14][7] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\uart_inst.fifo_rx_inst.mem[8][5] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\uart_inst.fifo_rx_inst.mem[12][7] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\uart_inst.fifo_tx_inst.mem[6][2] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\uart_inst.fifo_rx_inst.mem[0][5] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\uart_inst.fifo_rx_inst.mem[6][5] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\uart_inst.fifo_rx_inst.mem[0][6] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\uart_inst.fifo_rx_inst.mem[6][2] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\uart_inst.fifo_rx_inst.mem[8][6] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\uart_inst.fifo_rx_inst.mem[10][7] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\uart_inst.fifo_rx_inst.mem[10][0] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\uart_inst.fifo_rx_inst.mem[4][0] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\uart_inst.fifo_rx_inst.mem[8][3] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\uart_inst.fifo_rx_inst.mem[10][4] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\uart_inst.fifo_rx_inst.mem[2][7] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\uart_inst.fifo_rx_inst.mem[12][3] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\uart_inst.fifo_rx_inst.mem[14][0] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\uart_inst.fifo_rx_inst.mem[5][6] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\uart_inst.fifo_rx_inst.mem[0][3] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\uart_inst.fifo_rx_inst.mem[5][3] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\uart_inst.fifo_rx_inst.mem[2][0] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\uart_inst.fifo_rx_inst.mem[2][6] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\uart_inst.fifo_tx_inst.mem[6][4] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\uart_inst.fifo_rx_inst.mem[14][1] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\uart_inst.fifo_rx_inst.mem[12][1] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\uart_inst.fifo_rx_inst.mem[14][5] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\uart_inst.fifo_rx_inst.mem[10][5] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\uart_inst.fifo_rx_inst.mem[2][1] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\uart_inst.fifo_rx_inst.mem[5][5] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\uart_inst.fifo_tx_inst.mem[4][2] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\uart_inst.fifo_rx_inst.mem[0][1] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\uart_inst.fifo_rx_inst.mem[12][0] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\uart_inst.fifo_rx_inst.mem[1][6] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\uart_inst.fifo_rx_inst.mem[2][5] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\uart_inst.fifo_rx_inst.mem[1][5] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\uart_inst.fifo_tx_inst.mem[15][1] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\uart_inst.fifo_rx_inst.mem[14][4] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\uart_inst.fifo_rx_inst.mem[3][5] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\uart_inst.fifo_rx_inst.mem[1][3] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\uart_inst.fifo_rx_inst.mem[5][4] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\uart_inst.fifo_rx_inst.mem[6][4] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\uart_inst.fifo_rx_inst.mem[4][2] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\uart_inst.fifo_rx_inst.mem[12][2] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\uart_inst.fifo_tx_inst.mem[14][7] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\uart_inst.fifo_rx_inst.mem[3][6] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\uart_inst.fifo_rx_inst.mem[13][7] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\uart_inst.fifo_tx_inst.mem[4][4] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\uart_inst.fifo_tx_inst.mem[15][5] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\uart_inst.fifo_rx_inst.mem[5][7] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\uart_inst.fifo_rx_inst.mem[14][6] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\uart_inst.fifo_rx_inst.mem[12][6] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\uart_inst.fifo_rx_inst.mem[2][4] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\uart_inst.fifo_rx_inst.mem[1][2] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\uart_inst.fifo_rx_inst.mem[15][0] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[7] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0007_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\uart_inst.fifo_tx_inst.mem[14][6] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[5] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\uart_inst.fifo_rx_inst.mem[15][7] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\uart_inst.fifo_tx_inst.mem[12][5] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\uart_inst.fifo_tx_inst.mem[15][3] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\uart_inst.fifo_rx_inst.mem[5][0] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\uart_inst.fifo_rx_inst.mem[4][5] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\uart_inst.fifo_rx_inst.mem[12][4] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\uart_inst.fifo_rx_inst.mem[11][7] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\uart_inst.fifo_tx_inst.mem[14][5] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\uart_inst.uart_core_inst.uart_rx_inst.data_reg[2] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\uart_inst.fifo_rx_inst.mem[15][4] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\uart_inst.fifo_rx_inst.mem[5][1] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\uart_inst.uart_core_inst.uart_tx_inst.data_reg[6] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\uart_inst.fifo_tx_inst.mem[15][6] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\uart_inst.fifo_rx_inst.mem[3][3] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\uart_inst.fifo_rx_inst.mem[15][1] ),
    .X(net166));
 sky130_fd_sc_hd__buf_1 input1 (.A(PADDR[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(PWDATA[2]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(PWDATA[3]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(PWDATA[4]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(PWDATA[5]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(PWDATA[6]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(PWDATA[7]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(PWRITE),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(uart_rx),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(PADDR[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(PADDR[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(PADDR[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(PENABLE),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(PRESETn),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(PSEL),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(PWDATA[0]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(PWDATA[1]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_1039_),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(_1038_),
    .X(net376));
 sky130_fd_sc_hd__buf_1 max_cap27 (.A(_0706_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 max_cap28 (.A(_0616_),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 max_cap29 (.A(_0533_),
    .X(net29));
 sky130_fd_sc_hd__buf_4 max_cap30 (.A(_0524_),
    .X(net30));
 sky130_fd_sc_hd__buf_1 max_cap31 (.A(_0791_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 max_cap33 (.A(_0765_),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 max_cap34 (.A(_0590_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 max_cap35 (.A(_0406_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 max_cap36 (.A(_0864_),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 max_cap37 (.A(net375),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 max_cap38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 max_cap39 (.A(_1038_),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 max_cap40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 max_cap41 (.A(net377),
    .X(net41));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(PRDATA[0]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(PRDATA[1]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(PRDATA[2]));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(PRDATA[3]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(PRDATA[4]));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(PRDATA[5]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(PRDATA[6]));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net25),
    .X(PRDATA[7]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(uart_tx));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 uart_apb_wrapper_67 (.HI(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3 (.A(_0955_),
    .X(net377));
 sky130_fd_sc_hd__buf_1 wire32 (.A(_0765_),
    .X(net32));
 assign PRDATA[10] = net44;
 assign PRDATA[11] = net45;
 assign PRDATA[12] = net46;
 assign PRDATA[13] = net47;
 assign PRDATA[14] = net48;
 assign PRDATA[15] = net49;
 assign PRDATA[16] = net50;
 assign PRDATA[17] = net51;
 assign PRDATA[18] = net52;
 assign PRDATA[19] = net53;
 assign PRDATA[20] = net54;
 assign PRDATA[21] = net55;
 assign PRDATA[22] = net56;
 assign PRDATA[23] = net57;
 assign PRDATA[24] = net58;
 assign PRDATA[25] = net59;
 assign PRDATA[26] = net60;
 assign PRDATA[27] = net61;
 assign PRDATA[28] = net62;
 assign PRDATA[29] = net63;
 assign PRDATA[30] = net64;
 assign PRDATA[31] = net65;
 assign PRDATA[8] = net42;
 assign PRDATA[9] = net43;
 assign PREADY = net67;
 assign PSLVERR = net66;
endmodule

